
module system (
	clk_clk,
	reset_reset_n,
	vga_clk_clk,
	vga_reset_reset);	

	input		clk_clk;
	input		reset_reset_n;
	output		vga_clk_clk;
	output		vga_reset_reset;
endmodule
