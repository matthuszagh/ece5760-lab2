// system.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module system (
		input  wire  clk_clk,         //         clk.clk
		input  wire  reset_reset_n,   //       reset.reset_n
		output wire  vga_clk_ext_clk, // vga_clk_ext.clk
		output wire  vga_clk_int_clk  // vga_clk_int.clk
	);

	system_pll_0 pll_0 (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (vga_clk_int_clk), // outclk0.clk
		.outclk_1 (vga_clk_ext_clk), // outclk1.clk
		.locked   ()                 // (terminated)
	);

endmodule
