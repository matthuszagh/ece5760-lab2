// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition"

// DATE "05/18/2018 14:43:58"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module system (
	clk_clk,
	hps_io_hps_io_emac1_inst_TX_CLK,
	hps_io_hps_io_emac1_inst_TXD0,
	hps_io_hps_io_emac1_inst_TXD1,
	hps_io_hps_io_emac1_inst_TXD2,
	hps_io_hps_io_emac1_inst_TXD3,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_MDIO,
	hps_io_hps_io_emac1_inst_MDC,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_emac1_inst_TX_CTL,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_qspi_inst_IO0,
	hps_io_hps_io_qspi_inst_IO1,
	hps_io_hps_io_qspi_inst_IO2,
	hps_io_hps_io_qspi_inst_IO3,
	hps_io_hps_io_qspi_inst_SS0,
	hps_io_hps_io_qspi_inst_CLK,
	hps_io_hps_io_sdio_inst_CMD,
	hps_io_hps_io_sdio_inst_D0,
	hps_io_hps_io_sdio_inst_D1,
	hps_io_hps_io_sdio_inst_CLK,
	hps_io_hps_io_sdio_inst_D2,
	hps_io_hps_io_sdio_inst_D3,
	hps_io_hps_io_usb1_inst_D0,
	hps_io_hps_io_usb1_inst_D1,
	hps_io_hps_io_usb1_inst_D2,
	hps_io_hps_io_usb1_inst_D3,
	hps_io_hps_io_usb1_inst_D4,
	hps_io_hps_io_usb1_inst_D5,
	hps_io_hps_io_usb1_inst_D6,
	hps_io_hps_io_usb1_inst_D7,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_STP,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	hps_io_hps_io_spim1_inst_CLK,
	hps_io_hps_io_spim1_inst_MOSI,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_spim1_inst_SS0,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_uart0_inst_TX,
	hps_io_hps_io_i2c0_inst_SDA,
	hps_io_hps_io_i2c0_inst_SCL,
	hps_io_hps_io_i2c1_inst_SDA,
	hps_io_hps_io_i2c1_inst_SCL,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	ram_conduit_address,
	ram_conduit_chipselect,
	ram_conduit_clken,
	ram_conduit_write,
	ram_conduit_readdata,
	ram_conduit_writedata,
	ram_conduit_byteenable,
	reset_reset_n,
	vga_clk_ext_clk,
	vga_clk_int_clk)/* synthesis synthesis_greybox=0 */;
input 	clk_clk;
output 	hps_io_hps_io_emac1_inst_TX_CLK;
output 	hps_io_hps_io_emac1_inst_TXD0;
output 	hps_io_hps_io_emac1_inst_TXD1;
output 	hps_io_hps_io_emac1_inst_TXD2;
output 	hps_io_hps_io_emac1_inst_TXD3;
input 	hps_io_hps_io_emac1_inst_RXD0;
inout 	hps_io_hps_io_emac1_inst_MDIO;
output 	hps_io_hps_io_emac1_inst_MDC;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
output 	hps_io_hps_io_emac1_inst_TX_CTL;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
inout 	hps_io_hps_io_qspi_inst_IO0;
inout 	hps_io_hps_io_qspi_inst_IO1;
inout 	hps_io_hps_io_qspi_inst_IO2;
inout 	hps_io_hps_io_qspi_inst_IO3;
output 	hps_io_hps_io_qspi_inst_SS0;
output 	hps_io_hps_io_qspi_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_CMD;
inout 	hps_io_hps_io_sdio_inst_D0;
inout 	hps_io_hps_io_sdio_inst_D1;
output 	hps_io_hps_io_sdio_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_D2;
inout 	hps_io_hps_io_sdio_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D0;
inout 	hps_io_hps_io_usb1_inst_D1;
inout 	hps_io_hps_io_usb1_inst_D2;
inout 	hps_io_hps_io_usb1_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D4;
inout 	hps_io_hps_io_usb1_inst_D5;
inout 	hps_io_hps_io_usb1_inst_D6;
inout 	hps_io_hps_io_usb1_inst_D7;
input 	hps_io_hps_io_usb1_inst_CLK;
output 	hps_io_hps_io_usb1_inst_STP;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
output 	hps_io_hps_io_spim1_inst_CLK;
output 	hps_io_hps_io_spim1_inst_MOSI;
input 	hps_io_hps_io_spim1_inst_MISO;
output 	hps_io_hps_io_spim1_inst_SS0;
input 	hps_io_hps_io_uart0_inst_RX;
output 	hps_io_hps_io_uart0_inst_TX;
inout 	hps_io_hps_io_i2c0_inst_SDA;
inout 	hps_io_hps_io_i2c0_inst_SCL;
inout 	hps_io_hps_io_i2c1_inst_SDA;
inout 	hps_io_hps_io_i2c1_inst_SCL;
output 	[14:0] memory_mem_a;
output 	[2:0] memory_mem_ba;
output 	memory_mem_ck;
output 	memory_mem_ck_n;
output 	memory_mem_cke;
output 	memory_mem_cs_n;
output 	memory_mem_ras_n;
output 	memory_mem_cas_n;
output 	memory_mem_we_n;
output 	memory_mem_reset_n;
inout 	[31:0] memory_mem_dq;
inout 	[3:0] memory_mem_dqs;
inout 	[3:0] memory_mem_dqs_n;
output 	memory_mem_odt;
output 	[3:0] memory_mem_dm;
input 	memory_oct_rzqin;
input 	[3:0] ram_conduit_address;
input 	ram_conduit_chipselect;
input 	ram_conduit_clken;
input 	ram_conduit_write;
output 	[15:0] ram_conduit_readdata;
input 	[15:0] ram_conduit_writedata;
input 	[1:0] ram_conduit_byteenable;
input 	reset_reset_n;
output 	vga_clk_ext_clk;
output 	vga_clk_int_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_0|fpga_interfaces|h2f_rst_n[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_BREADY[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_RREADY[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WLAST[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARBURST[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARBURST[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARSIZE[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARSIZE[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARSIZE[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWBURST[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWBURST[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWSIZE[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWSIZE[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWSIZE[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[12] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[13] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[14] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[15] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[16] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[17] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[18] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[19] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[20] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[21] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[22] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[23] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[24] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[25] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[26] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[27] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[28] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[29] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[30] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[31] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[3] ;
wire \ram|the_altsyncram|auto_generated|q_a[0] ;
wire \ram|the_altsyncram|auto_generated|q_b[0] ;
wire \ram|the_altsyncram|auto_generated|q_a[1] ;
wire \ram|the_altsyncram|auto_generated|q_b[1] ;
wire \ram|the_altsyncram|auto_generated|q_a[2] ;
wire \ram|the_altsyncram|auto_generated|q_b[2] ;
wire \ram|the_altsyncram|auto_generated|q_a[3] ;
wire \ram|the_altsyncram|auto_generated|q_b[3] ;
wire \ram|the_altsyncram|auto_generated|q_a[4] ;
wire \ram|the_altsyncram|auto_generated|q_b[4] ;
wire \ram|the_altsyncram|auto_generated|q_a[5] ;
wire \ram|the_altsyncram|auto_generated|q_b[5] ;
wire \ram|the_altsyncram|auto_generated|q_a[6] ;
wire \ram|the_altsyncram|auto_generated|q_b[6] ;
wire \ram|the_altsyncram|auto_generated|q_a[7] ;
wire \ram|the_altsyncram|auto_generated|q_b[7] ;
wire \ram|the_altsyncram|auto_generated|q_a[8] ;
wire \ram|the_altsyncram|auto_generated|q_b[8] ;
wire \ram|the_altsyncram|auto_generated|q_a[9] ;
wire \ram|the_altsyncram|auto_generated|q_b[9] ;
wire \ram|the_altsyncram|auto_generated|q_a[10] ;
wire \ram|the_altsyncram|auto_generated|q_b[10] ;
wire \ram|the_altsyncram|auto_generated|q_a[11] ;
wire \ram|the_altsyncram|auto_generated|q_b[11] ;
wire \ram|the_altsyncram|auto_generated|q_a[12] ;
wire \ram|the_altsyncram|auto_generated|q_b[12] ;
wire \ram|the_altsyncram|auto_generated|q_a[13] ;
wire \ram|the_altsyncram|auto_generated|q_b[13] ;
wire \ram|the_altsyncram|auto_generated|q_a[14] ;
wire \ram|the_altsyncram|auto_generated|q_b[14] ;
wire \ram|the_altsyncram|auto_generated|q_a[15] ;
wire \ram|the_altsyncram|auto_generated|q_b[15] ;
wire \pll_0|altera_pll_i|outclk_wire[1] ;
wire \pll_0|altera_pll_i|outclk_wire[0] ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[1]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|cmd_mux|sink1_ready~combout ;
wire \mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|awready~0_combout ;
wire \mm_interconnect_0|rsp_demux|src0_valid~1_combout ;
wire \mm_interconnect_0|ram_s1_agent|uncompressor|source_endofpacket~combout ;
wire \mm_interconnect_0|rsp_demux|src1_valid~0_combout ;
wire \mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|wready~0_combout ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][70]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][71]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][72]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][73]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][79]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][80]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][81]~q ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[0]~0_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[1]~1_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[2]~2_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[3]~3_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[4]~4_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[5]~5_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[6]~6_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[7]~7_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[8]~8_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[9]~9_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[10]~10_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[11]~11_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[12]~12_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[13]~13_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[14]~14_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[15]~15_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~16_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~17_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~18_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~19_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~20_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~21_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~22_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~23_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~24_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~25_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~26_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~27_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~28_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~29_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~30_combout ;
wire \mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~31_combout ;
wire \mm_interconnect_0|ram_s1_agent|m0_write~1_combout ;
wire \rst_controller_001|r_early_rst~q ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[16]~0_combout ;
wire \mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[17]~1_combout ;
wire \rst_controller|merged_reset~0_combout ;
wire \rst_controller_001|r_sync_rst~q ;
wire \rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \~GND~combout ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;
wire \hps_0|hps_io|border|intermediate[0] ;
wire \hps_0|hps_io|border|intermediate[1] ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;
wire \hps_0|hps_io|border|emac1_inst~emac_phy_txd ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;
wire \hps_0|hps_io|border|qspi_inst~O_QSPI_SCLK ;
wire \hps_0|hps_io|border|intermediate[2] ;
wire \hps_0|hps_io|border|intermediate[4] ;
wire \hps_0|hps_io|border|intermediate[6] ;
wire \hps_0|hps_io|border|intermediate[8] ;
wire \hps_0|hps_io|border|intermediate[3] ;
wire \hps_0|hps_io|border|intermediate[5] ;
wire \hps_0|hps_io|border|intermediate[7] ;
wire \hps_0|hps_io|border|intermediate[9] ;
wire \hps_0|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;
wire \hps_0|hps_io|border|sdio_inst~sdmmc_cclk ;
wire \hps_0|hps_io|border|intermediate[10] ;
wire \hps_0|hps_io|border|intermediate[11] ;
wire \hps_0|hps_io|border|intermediate[12] ;
wire \hps_0|hps_io|border|intermediate[14] ;
wire \hps_0|hps_io|border|intermediate[16] ;
wire \hps_0|hps_io|border|intermediate[18] ;
wire \hps_0|hps_io|border|intermediate[13] ;
wire \hps_0|hps_io|border|intermediate[15] ;
wire \hps_0|hps_io|border|intermediate[17] ;
wire \hps_0|hps_io|border|intermediate[19] ;
wire \hps_0|hps_io|border|usb1_inst~usb_ulpi_stp ;
wire \hps_0|hps_io|border|intermediate[20] ;
wire \hps_0|hps_io|border|intermediate[22] ;
wire \hps_0|hps_io|border|intermediate[24] ;
wire \hps_0|hps_io|border|intermediate[26] ;
wire \hps_0|hps_io|border|intermediate[28] ;
wire \hps_0|hps_io|border|intermediate[30] ;
wire \hps_0|hps_io|border|intermediate[32] ;
wire \hps_0|hps_io|border|intermediate[34] ;
wire \hps_0|hps_io|border|intermediate[21] ;
wire \hps_0|hps_io|border|intermediate[23] ;
wire \hps_0|hps_io|border|intermediate[25] ;
wire \hps_0|hps_io|border|intermediate[27] ;
wire \hps_0|hps_io|border|intermediate[29] ;
wire \hps_0|hps_io|border|intermediate[31] ;
wire \hps_0|hps_io|border|intermediate[33] ;
wire \hps_0|hps_io|border|intermediate[35] ;
wire \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;
wire \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;
wire \hps_0|hps_io|border|intermediate[36] ;
wire \hps_0|hps_io|border|intermediate[37] ;
wire \hps_0|hps_io|border|uart0_inst~uart_txd ;
wire \hps_0|hps_io|border|intermediate[39] ;
wire \hps_0|hps_io|border|intermediate[38] ;
wire \hps_0|hps_io|border|intermediate[41] ;
wire \hps_0|hps_io|border|intermediate[40] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o ;
wire \clk_clk~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD0~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD1~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD2~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD3~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CLK~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CTL~input_o ;
wire \hps_io_hps_io_spim1_inst_MISO~input_o ;
wire \hps_io_hps_io_uart0_inst_RX~input_o ;
wire \hps_io_hps_io_usb1_inst_CLK~input_o ;
wire \hps_io_hps_io_usb1_inst_DIR~input_o ;
wire \hps_io_hps_io_usb1_inst_NXT~input_o ;
wire \memory_oct_rzqin~input_o ;
wire \ram_conduit_chipselect~input_o ;
wire \ram_conduit_write~input_o ;
wire \ram_conduit_clken~input_o ;
wire \ram_conduit_writedata[0]~input_o ;
wire \ram_conduit_address[0]~input_o ;
wire \ram_conduit_address[1]~input_o ;
wire \ram_conduit_address[2]~input_o ;
wire \ram_conduit_address[3]~input_o ;
wire \ram_conduit_byteenable[0]~input_o ;
wire \ram_conduit_writedata[1]~input_o ;
wire \ram_conduit_writedata[2]~input_o ;
wire \ram_conduit_writedata[3]~input_o ;
wire \ram_conduit_writedata[4]~input_o ;
wire \ram_conduit_writedata[5]~input_o ;
wire \ram_conduit_writedata[6]~input_o ;
wire \ram_conduit_writedata[7]~input_o ;
wire \ram_conduit_writedata[8]~input_o ;
wire \ram_conduit_byteenable[1]~input_o ;
wire \ram_conduit_writedata[9]~input_o ;
wire \ram_conduit_writedata[10]~input_o ;
wire \ram_conduit_writedata[11]~input_o ;
wire \ram_conduit_writedata[12]~input_o ;
wire \ram_conduit_writedata[13]~input_o ;
wire \ram_conduit_writedata[14]~input_o ;
wire \ram_conduit_writedata[15]~input_o ;
wire \reset_reset_n~input_o ;


system_system_mm_interconnect_0 mm_interconnect_0(
	.h2f_lw_ARVALID_0(\hps_0|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\hps_0|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\hps_0|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\hps_0|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\hps_0|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\hps_0|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\hps_0|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\hps_0|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\hps_0|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\hps_0|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\hps_0|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARBURST_0(\hps_0|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\hps_0|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\hps_0|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\hps_0|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\hps_0|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\hps_0|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\hps_0|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\hps_0|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\hps_0|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\hps_0|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\hps_0|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\hps_0|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\hps_0|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\hps_0|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\hps_0|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\hps_0|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\hps_0|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\hps_0|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\hps_0|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\hps_0|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\hps_0|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\hps_0|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\hps_0|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWBURST_0(\hps_0|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\hps_0|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\hps_0|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\hps_0|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\hps_0|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\hps_0|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\hps_0|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\hps_0|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\hps_0|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\hps_0|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\hps_0|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\hps_0|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\hps_0|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\hps_0|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\hps_0|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\hps_0|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\hps_0|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\hps_0|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\hps_0|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\hps_0|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\hps_0|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\hps_0|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\hps_0|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\hps_0|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\hps_0|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\hps_0|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\hps_0|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\hps_0|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\hps_0|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\hps_0|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\hps_0|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\hps_0|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\hps_0|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\hps_0|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\hps_0|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\hps_0|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\hps_0|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\hps_0|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\hps_0|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\hps_0|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\hps_0|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\hps_0|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\hps_0|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\hps_0|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\hps_0|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\hps_0|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\hps_0|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\hps_0|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\hps_0|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\hps_0|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\hps_0|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\hps_0|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\hps_0|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\hps_0|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.q_a_0(\ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_8(\ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_10(\ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_11(\ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_12(\ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\ram|the_altsyncram|auto_generated|q_a[15] ),
	.in_data_reg_0(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_1(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[1]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.in_data_reg_1(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.sink1_ready(\mm_interconnect_0|cmd_mux|sink1_ready~combout ),
	.hps_0_h2f_lw_axi_master_awready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|awready~0_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux|src0_valid~1_combout ),
	.source_endofpacket(\mm_interconnect_0|ram_s1_agent|uncompressor|source_endofpacket~combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux|src1_valid~0_combout ),
	.hps_0_h2f_lw_axi_master_wready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|wready~0_combout ),
	.mem_70_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][70]~q ),
	.mem_71_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][71]~q ),
	.mem_72_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][72]~q ),
	.mem_73_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][73]~q ),
	.mem_74_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_75_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_76_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_77_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_78_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_79_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][79]~q ),
	.mem_80_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][80]~q ),
	.mem_81_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][81]~q ),
	.out_data_0(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[0]~0_combout ),
	.out_data_1(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[1]~1_combout ),
	.out_data_2(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[2]~2_combout ),
	.out_data_3(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[3]~3_combout ),
	.out_data_4(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[4]~4_combout ),
	.out_data_5(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[5]~5_combout ),
	.out_data_6(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[6]~6_combout ),
	.out_data_7(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[7]~7_combout ),
	.out_data_8(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[8]~8_combout ),
	.out_data_9(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[9]~9_combout ),
	.out_data_10(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[10]~10_combout ),
	.out_data_11(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[11]~11_combout ),
	.out_data_12(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[12]~12_combout ),
	.out_data_13(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[13]~13_combout ),
	.out_data_14(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[14]~14_combout ),
	.out_data_15(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[15]~15_combout ),
	.ShiftLeft2(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~16_combout ),
	.ShiftLeft21(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~17_combout ),
	.ShiftLeft22(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~18_combout ),
	.ShiftLeft23(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~19_combout ),
	.ShiftLeft24(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~20_combout ),
	.ShiftLeft25(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~21_combout ),
	.ShiftLeft26(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~22_combout ),
	.ShiftLeft27(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~23_combout ),
	.ShiftLeft28(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~24_combout ),
	.ShiftLeft29(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~25_combout ),
	.ShiftLeft210(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~26_combout ),
	.ShiftLeft211(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~27_combout ),
	.ShiftLeft212(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~28_combout ),
	.ShiftLeft213(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~29_combout ),
	.ShiftLeft214(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~30_combout ),
	.ShiftLeft215(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~31_combout ),
	.m0_write(\mm_interconnect_0|ram_s1_agent|m0_write~1_combout ),
	.source0_data_16(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[16]~0_combout ),
	.source0_data_17(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[17]~1_combout ),
	.r_sync_rst(\rst_controller_001|r_sync_rst~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

system_system_ram ram(
	.q_a_0(\ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_b_0(\ram|the_altsyncram|auto_generated|q_b[0] ),
	.q_a_1(\ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_b_1(\ram|the_altsyncram|auto_generated|q_b[1] ),
	.q_a_2(\ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_b_2(\ram|the_altsyncram|auto_generated|q_b[2] ),
	.q_a_3(\ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_b_3(\ram|the_altsyncram|auto_generated|q_b[3] ),
	.q_a_4(\ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_b_4(\ram|the_altsyncram|auto_generated|q_b[4] ),
	.q_a_5(\ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_b_5(\ram|the_altsyncram|auto_generated|q_b[5] ),
	.q_a_6(\ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_b_6(\ram|the_altsyncram|auto_generated|q_b[6] ),
	.q_a_7(\ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_b_7(\ram|the_altsyncram|auto_generated|q_b[7] ),
	.q_a_8(\ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_b_8(\ram|the_altsyncram|auto_generated|q_b[8] ),
	.q_a_9(\ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_b_9(\ram|the_altsyncram|auto_generated|q_b[9] ),
	.q_a_10(\ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_b_10(\ram|the_altsyncram|auto_generated|q_b[10] ),
	.q_a_11(\ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_b_11(\ram|the_altsyncram|auto_generated|q_b[11] ),
	.q_a_12(\ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_b_12(\ram|the_altsyncram|auto_generated|q_b[12] ),
	.q_a_13(\ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_b_13(\ram|the_altsyncram|auto_generated|q_b[13] ),
	.q_a_14(\ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_b_14(\ram|the_altsyncram|auto_generated|q_b[14] ),
	.q_a_15(\ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_b_15(\ram|the_altsyncram|auto_generated|q_b[15] ),
	.in_data_reg_0(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_1(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[1]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.in_data_reg_1(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.m0_write(\mm_interconnect_0|ram_s1_agent|m0_write~1_combout ),
	.r_early_rst(\rst_controller_001|r_early_rst~q ),
	.source0_data_16(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[16]~0_combout ),
	.source0_data_17(\mm_interconnect_0|ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[17]~1_combout ),
	.clk_clk(\clk_clk~input_o ),
	.ram_conduit_chipselect(\ram_conduit_chipselect~input_o ),
	.ram_conduit_write(\ram_conduit_write~input_o ),
	.ram_conduit_clken(\ram_conduit_clken~input_o ),
	.ram_conduit_writedata_0(\ram_conduit_writedata[0]~input_o ),
	.ram_conduit_address_0(\ram_conduit_address[0]~input_o ),
	.ram_conduit_address_1(\ram_conduit_address[1]~input_o ),
	.ram_conduit_address_2(\ram_conduit_address[2]~input_o ),
	.ram_conduit_address_3(\ram_conduit_address[3]~input_o ),
	.ram_conduit_byteenable_0(\ram_conduit_byteenable[0]~input_o ),
	.ram_conduit_writedata_1(\ram_conduit_writedata[1]~input_o ),
	.ram_conduit_writedata_2(\ram_conduit_writedata[2]~input_o ),
	.ram_conduit_writedata_3(\ram_conduit_writedata[3]~input_o ),
	.ram_conduit_writedata_4(\ram_conduit_writedata[4]~input_o ),
	.ram_conduit_writedata_5(\ram_conduit_writedata[5]~input_o ),
	.ram_conduit_writedata_6(\ram_conduit_writedata[6]~input_o ),
	.ram_conduit_writedata_7(\ram_conduit_writedata[7]~input_o ),
	.ram_conduit_writedata_8(\ram_conduit_writedata[8]~input_o ),
	.ram_conduit_byteenable_1(\ram_conduit_byteenable[1]~input_o ),
	.ram_conduit_writedata_9(\ram_conduit_writedata[9]~input_o ),
	.ram_conduit_writedata_10(\ram_conduit_writedata[10]~input_o ),
	.ram_conduit_writedata_11(\ram_conduit_writedata[11]~input_o ),
	.ram_conduit_writedata_12(\ram_conduit_writedata[12]~input_o ),
	.ram_conduit_writedata_13(\ram_conduit_writedata[13]~input_o ),
	.ram_conduit_writedata_14(\ram_conduit_writedata[14]~input_o ),
	.ram_conduit_writedata_15(\ram_conduit_writedata[15]~input_o ));

system_system_pll_0 pll_0(
	.outclk_wire_1(\pll_0|altera_pll_i|outclk_wire[1] ),
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.merged_reset(\rst_controller|merged_reset~0_combout ),
	.clk_clk(\clk_clk~input_o ));

system_altera_reset_controller_2 rst_controller_002(
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ));

system_altera_reset_controller_1 rst_controller_001(
	.r_early_rst1(\rst_controller_001|r_early_rst~q ),
	.merged_reset(\rst_controller|merged_reset~0_combout ),
	.r_sync_rst1(\rst_controller_001|r_sync_rst~q ),
	.clk_clk(\clk_clk~input_o ));

system_altera_reset_controller rst_controller(
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.merged_reset(\rst_controller|merged_reset~0_combout ),
	.reset_reset_n(\reset_reset_n~input_o ));

system_system_hps_0 hps_0(
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.h2f_lw_ARVALID_0(\hps_0|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\hps_0|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\hps_0|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\hps_0|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\hps_0|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\hps_0|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\hps_0|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\hps_0|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\hps_0|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\hps_0|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\hps_0|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARBURST_0(\hps_0|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\hps_0|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\hps_0|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\hps_0|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\hps_0|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\hps_0|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\hps_0|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\hps_0|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\hps_0|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\hps_0|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\hps_0|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\hps_0|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\hps_0|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\hps_0|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\hps_0|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\hps_0|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\hps_0|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\hps_0|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\hps_0|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\hps_0|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\hps_0|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\hps_0|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\hps_0|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWBURST_0(\hps_0|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\hps_0|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\hps_0|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\hps_0|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\hps_0|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\hps_0|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\hps_0|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\hps_0|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\hps_0|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\hps_0|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\hps_0|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\hps_0|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\hps_0|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\hps_0|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\hps_0|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\hps_0|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\hps_0|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\hps_0|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\hps_0|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\hps_0|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\hps_0|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\hps_0|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\hps_0|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\hps_0|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\hps_0|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\hps_0|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\hps_0|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\hps_0|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\hps_0|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\hps_0|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\hps_0|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\hps_0|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\hps_0|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\hps_0|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\hps_0|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\hps_0|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\hps_0|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\hps_0|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\hps_0|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\hps_0|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\hps_0|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\hps_0|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\hps_0|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\hps_0|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\hps_0|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\hps_0|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\hps_0|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\hps_0|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\hps_0|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\hps_0|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\hps_0|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\hps_0|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\hps_0|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\hps_0|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.sink1_ready(\mm_interconnect_0|cmd_mux|sink1_ready~combout ),
	.awready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|awready~0_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux|src0_valid~1_combout ),
	.source_endofpacket(\mm_interconnect_0|ram_s1_agent|uncompressor|source_endofpacket~combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux|src1_valid~0_combout ),
	.wready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|wready~0_combout ),
	.mem_70_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][70]~q ),
	.mem_71_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][71]~q ),
	.mem_72_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][72]~q ),
	.mem_73_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][73]~q ),
	.mem_74_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_75_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_76_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_77_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_78_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_79_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][79]~q ),
	.mem_80_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][80]~q ),
	.mem_81_0(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem[0][81]~q ),
	.out_data_0(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[0]~0_combout ),
	.out_data_1(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[1]~1_combout ),
	.out_data_2(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[2]~2_combout ),
	.out_data_3(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[3]~3_combout ),
	.out_data_4(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[4]~4_combout ),
	.out_data_5(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[5]~5_combout ),
	.out_data_6(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[6]~6_combout ),
	.out_data_7(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[7]~7_combout ),
	.out_data_8(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[8]~8_combout ),
	.out_data_9(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[9]~9_combout ),
	.out_data_10(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[10]~10_combout ),
	.out_data_11(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[11]~11_combout ),
	.out_data_12(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[12]~12_combout ),
	.out_data_13(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[13]~13_combout ),
	.out_data_14(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[14]~14_combout ),
	.out_data_15(\mm_interconnect_0|ram_s1_rsp_width_adapter|out_data[15]~15_combout ),
	.ShiftLeft2(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~16_combout ),
	.ShiftLeft21(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~17_combout ),
	.ShiftLeft22(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~18_combout ),
	.ShiftLeft23(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~19_combout ),
	.ShiftLeft24(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~20_combout ),
	.ShiftLeft25(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~21_combout ),
	.ShiftLeft26(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~22_combout ),
	.ShiftLeft27(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~23_combout ),
	.ShiftLeft28(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~24_combout ),
	.ShiftLeft29(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~25_combout ),
	.ShiftLeft210(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~26_combout ),
	.ShiftLeft211(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~27_combout ),
	.ShiftLeft212(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~28_combout ),
	.ShiftLeft213(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~29_combout ),
	.ShiftLeft214(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~30_combout ),
	.ShiftLeft215(\mm_interconnect_0|ram_s1_rsp_width_adapter|ShiftLeft2~31_combout ),
	.emac1_inst(\hps_0|hps_io|border|emac1_inst~O_EMAC_CLK_TX ),
	.emac1_inst1(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ),
	.intermediate_0(\hps_0|hps_io|border|intermediate[0] ),
	.intermediate_1(\hps_0|hps_io|border|intermediate[1] ),
	.emac1_inst2(\hps_0|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ),
	.emac1_inst3(\hps_0|hps_io|border|emac1_inst~emac_phy_txd ),
	.emac1_inst4(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ),
	.emac1_inst5(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ),
	.emac1_inst6(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ),
	.qspi_inst(\hps_0|hps_io|border|qspi_inst~O_QSPI_SCLK ),
	.intermediate_2(\hps_0|hps_io|border|intermediate[2] ),
	.intermediate_4(\hps_0|hps_io|border|intermediate[4] ),
	.intermediate_6(\hps_0|hps_io|border|intermediate[6] ),
	.intermediate_8(\hps_0|hps_io|border|intermediate[8] ),
	.intermediate_3(\hps_0|hps_io|border|intermediate[3] ),
	.intermediate_5(\hps_0|hps_io|border|intermediate[5] ),
	.intermediate_7(\hps_0|hps_io|border|intermediate[7] ),
	.intermediate_9(\hps_0|hps_io|border|intermediate[9] ),
	.qspi_inst1(\hps_0|hps_io|border|qspi_inst~O_QSPI_SS_N0 ),
	.sdio_inst(\hps_0|hps_io|border|sdio_inst~sdmmc_cclk ),
	.intermediate_10(\hps_0|hps_io|border|intermediate[10] ),
	.intermediate_11(\hps_0|hps_io|border|intermediate[11] ),
	.intermediate_12(\hps_0|hps_io|border|intermediate[12] ),
	.intermediate_14(\hps_0|hps_io|border|intermediate[14] ),
	.intermediate_16(\hps_0|hps_io|border|intermediate[16] ),
	.intermediate_18(\hps_0|hps_io|border|intermediate[18] ),
	.intermediate_13(\hps_0|hps_io|border|intermediate[13] ),
	.intermediate_15(\hps_0|hps_io|border|intermediate[15] ),
	.intermediate_17(\hps_0|hps_io|border|intermediate[17] ),
	.intermediate_19(\hps_0|hps_io|border|intermediate[19] ),
	.usb1_inst(\hps_0|hps_io|border|usb1_inst~usb_ulpi_stp ),
	.intermediate_20(\hps_0|hps_io|border|intermediate[20] ),
	.intermediate_22(\hps_0|hps_io|border|intermediate[22] ),
	.intermediate_24(\hps_0|hps_io|border|intermediate[24] ),
	.intermediate_26(\hps_0|hps_io|border|intermediate[26] ),
	.intermediate_28(\hps_0|hps_io|border|intermediate[28] ),
	.intermediate_30(\hps_0|hps_io|border|intermediate[30] ),
	.intermediate_32(\hps_0|hps_io|border|intermediate[32] ),
	.intermediate_34(\hps_0|hps_io|border|intermediate[34] ),
	.intermediate_21(\hps_0|hps_io|border|intermediate[21] ),
	.intermediate_23(\hps_0|hps_io|border|intermediate[23] ),
	.intermediate_25(\hps_0|hps_io|border|intermediate[25] ),
	.intermediate_27(\hps_0|hps_io|border|intermediate[27] ),
	.intermediate_29(\hps_0|hps_io|border|intermediate[29] ),
	.intermediate_31(\hps_0|hps_io|border|intermediate[31] ),
	.intermediate_33(\hps_0|hps_io|border|intermediate[33] ),
	.intermediate_35(\hps_0|hps_io|border|intermediate[35] ),
	.spim1_inst(\hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ),
	.spim1_inst1(\hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ),
	.intermediate_36(\hps_0|hps_io|border|intermediate[36] ),
	.intermediate_37(\hps_0|hps_io|border|intermediate[37] ),
	.uart0_inst(\hps_0|hps_io|border|uart0_inst~uart_txd ),
	.intermediate_39(\hps_0|hps_io|border|intermediate[39] ),
	.intermediate_38(\hps_0|hps_io|border|intermediate[38] ),
	.intermediate_41(\hps_0|hps_io|border|intermediate[41] ),
	.intermediate_40(\hps_0|hps_io|border|intermediate[40] ),
	.parallelterminationcontrol_0(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ),
	.parallelterminationcontrol_1(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ),
	.parallelterminationcontrol_2(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ),
	.parallelterminationcontrol_3(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ),
	.parallelterminationcontrol_4(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ),
	.parallelterminationcontrol_5(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ),
	.parallelterminationcontrol_6(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ),
	.parallelterminationcontrol_7(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ),
	.parallelterminationcontrol_8(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ),
	.parallelterminationcontrol_9(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ),
	.parallelterminationcontrol_10(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ),
	.parallelterminationcontrol_11(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ),
	.parallelterminationcontrol_12(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ),
	.parallelterminationcontrol_13(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ),
	.parallelterminationcontrol_14(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ),
	.parallelterminationcontrol_15(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ),
	.seriesterminationcontrol_0(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ),
	.seriesterminationcontrol_1(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ),
	.seriesterminationcontrol_2(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ),
	.seriesterminationcontrol_3(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ),
	.seriesterminationcontrol_4(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ),
	.seriesterminationcontrol_5(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ),
	.seriesterminationcontrol_6(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ),
	.seriesterminationcontrol_7(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ),
	.seriesterminationcontrol_8(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ),
	.seriesterminationcontrol_9(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ),
	.seriesterminationcontrol_10(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ),
	.seriesterminationcontrol_11(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ),
	.seriesterminationcontrol_12(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ),
	.seriesterminationcontrol_13(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ),
	.seriesterminationcontrol_14(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ),
	.seriesterminationcontrol_15(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ),
	.dqsin(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dataout_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ),
	.dataout_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ),
	.dataout_2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ),
	.dataout_3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ),
	.dataout_4(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ),
	.dataout_5(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ),
	.dataout_6(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ),
	.dataout_7(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ),
	.dataout_8(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ),
	.dataout_9(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ),
	.dataout_10(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ),
	.dataout_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ),
	.dataout_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ),
	.dataout_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ),
	.dataout_14(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ),
	.dataout_01(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ),
	.dataout_15(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ),
	.dataout_21(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ),
	.dataout_16(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ),
	.dataout_02(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ),
	.dataout_31(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ),
	.dataout_41(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ),
	.dataout_51(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ),
	.dataout_03(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ),
	.dataout_22(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ),
	.extra_output_pad_gen0delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.wire_pseudo_diffa_o_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.wire_pseudo_diffa_obar_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.wire_pseudo_diffa_oeout_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.wire_pseudo_diffa_oebout_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.pad_gen0delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.os(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.hps_io_emac1_inst_MDIO_0(\hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ),
	.hps_io_qspi_inst_IO0_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ),
	.hps_io_qspi_inst_IO1_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ),
	.hps_io_qspi_inst_IO2_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ),
	.hps_io_qspi_inst_IO3_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ),
	.hps_io_sdio_inst_CMD_0(\hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ),
	.hps_io_sdio_inst_D0_0(\hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ),
	.hps_io_sdio_inst_D1_0(\hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ),
	.hps_io_sdio_inst_D2_0(\hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ),
	.hps_io_sdio_inst_D3_0(\hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D0_0(\hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ),
	.hps_io_usb1_inst_D1_0(\hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ),
	.hps_io_usb1_inst_D2_0(\hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ),
	.hps_io_usb1_inst_D3_0(\hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D4_0(\hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ),
	.hps_io_usb1_inst_D5_0(\hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ),
	.hps_io_usb1_inst_D6_0(\hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ),
	.hps_io_usb1_inst_D7_0(\hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ),
	.hps_io_i2c0_inst_SDA_0(\hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o ),
	.hps_io_i2c0_inst_SCL_0(\hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o ),
	.hps_io_i2c1_inst_SDA_0(\hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o ),
	.hps_io_i2c1_inst_SCL_0(\hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o ),
	.clk_clk(\clk_clk~input_o ),
	.hps_io_hps_io_emac1_inst_RXD0(\hps_io_hps_io_emac1_inst_RXD0~input_o ),
	.hps_io_hps_io_emac1_inst_RXD1(\hps_io_hps_io_emac1_inst_RXD1~input_o ),
	.hps_io_hps_io_emac1_inst_RXD2(\hps_io_hps_io_emac1_inst_RXD2~input_o ),
	.hps_io_hps_io_emac1_inst_RXD3(\hps_io_hps_io_emac1_inst_RXD3~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CLK(\hps_io_hps_io_emac1_inst_RX_CLK~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CTL(\hps_io_hps_io_emac1_inst_RX_CTL~input_o ),
	.hps_io_hps_io_spim1_inst_MISO(\hps_io_hps_io_spim1_inst_MISO~input_o ),
	.hps_io_hps_io_uart0_inst_RX(\hps_io_hps_io_uart0_inst_RX~input_o ),
	.hps_io_hps_io_usb1_inst_CLK(\hps_io_hps_io_usb1_inst_CLK~input_o ),
	.hps_io_hps_io_usb1_inst_DIR(\hps_io_hps_io_usb1_inst_DIR~input_o ),
	.hps_io_hps_io_usb1_inst_NXT(\hps_io_hps_io_usb1_inst_NXT~input_o ),
	.memory_oct_rzqin(\memory_oct_rzqin~input_o ));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[3]),
	.ibar(memory_mem_dqs_n[3]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[24]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[25]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[26]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[27]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[28]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[29]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[30]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[31]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[2]),
	.ibar(memory_mem_dqs_n[2]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[16]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[17]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[18]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[19]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[20]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[21]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[22]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[23]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[1]),
	.ibar(memory_mem_dqs_n[1]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[8]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[9]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[10]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[11]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[12]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[13]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[14]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[15]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[0]),
	.ibar(memory_mem_dqs_n[0]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[0]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[1]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[2]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[3]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[4]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[5]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[6]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[7]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

assign \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o  = hps_io_hps_io_emac1_inst_MDIO;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o  = hps_io_hps_io_qspi_inst_IO0;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o  = hps_io_hps_io_qspi_inst_IO1;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o  = hps_io_hps_io_qspi_inst_IO2;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o  = hps_io_hps_io_qspi_inst_IO3;

assign \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o  = hps_io_hps_io_sdio_inst_CMD;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~input_o  = hps_io_hps_io_sdio_inst_D0;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~input_o  = hps_io_hps_io_sdio_inst_D1;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~input_o  = hps_io_hps_io_sdio_inst_D2;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~input_o  = hps_io_hps_io_sdio_inst_D3;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~input_o  = hps_io_hps_io_usb1_inst_D0;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~input_o  = hps_io_hps_io_usb1_inst_D1;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~input_o  = hps_io_hps_io_usb1_inst_D2;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~input_o  = hps_io_hps_io_usb1_inst_D3;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~input_o  = hps_io_hps_io_usb1_inst_D4;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~input_o  = hps_io_hps_io_usb1_inst_D5;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~input_o  = hps_io_hps_io_usb1_inst_D6;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~input_o  = hps_io_hps_io_usb1_inst_D7;

assign \hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o  = hps_io_hps_io_i2c0_inst_SDA;

assign \hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o  = hps_io_hps_io_i2c0_inst_SCL;

assign \hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o  = hps_io_hps_io_i2c1_inst_SDA;

assign \hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o  = hps_io_hps_io_i2c1_inst_SCL;

assign \clk_clk~input_o  = clk_clk;

assign \hps_io_hps_io_emac1_inst_RXD0~input_o  = hps_io_hps_io_emac1_inst_RXD0;

assign \hps_io_hps_io_emac1_inst_RXD1~input_o  = hps_io_hps_io_emac1_inst_RXD1;

assign \hps_io_hps_io_emac1_inst_RXD2~input_o  = hps_io_hps_io_emac1_inst_RXD2;

assign \hps_io_hps_io_emac1_inst_RXD3~input_o  = hps_io_hps_io_emac1_inst_RXD3;

assign \hps_io_hps_io_emac1_inst_RX_CLK~input_o  = hps_io_hps_io_emac1_inst_RX_CLK;

assign \hps_io_hps_io_emac1_inst_RX_CTL~input_o  = hps_io_hps_io_emac1_inst_RX_CTL;

assign \hps_io_hps_io_spim1_inst_MISO~input_o  = hps_io_hps_io_spim1_inst_MISO;

assign \hps_io_hps_io_uart0_inst_RX~input_o  = hps_io_hps_io_uart0_inst_RX;

assign \hps_io_hps_io_usb1_inst_CLK~input_o  = hps_io_hps_io_usb1_inst_CLK;

assign \hps_io_hps_io_usb1_inst_DIR~input_o  = hps_io_hps_io_usb1_inst_DIR;

assign \hps_io_hps_io_usb1_inst_NXT~input_o  = hps_io_hps_io_usb1_inst_NXT;

assign \memory_oct_rzqin~input_o  = memory_oct_rzqin;

assign \ram_conduit_chipselect~input_o  = ram_conduit_chipselect;

assign \ram_conduit_write~input_o  = ram_conduit_write;

assign \ram_conduit_clken~input_o  = ram_conduit_clken;

assign \ram_conduit_writedata[0]~input_o  = ram_conduit_writedata[0];

assign \ram_conduit_address[0]~input_o  = ram_conduit_address[0];

assign \ram_conduit_address[1]~input_o  = ram_conduit_address[1];

assign \ram_conduit_address[2]~input_o  = ram_conduit_address[2];

assign \ram_conduit_address[3]~input_o  = ram_conduit_address[3];

assign \ram_conduit_byteenable[0]~input_o  = ram_conduit_byteenable[0];

assign \ram_conduit_writedata[1]~input_o  = ram_conduit_writedata[1];

assign \ram_conduit_writedata[2]~input_o  = ram_conduit_writedata[2];

assign \ram_conduit_writedata[3]~input_o  = ram_conduit_writedata[3];

assign \ram_conduit_writedata[4]~input_o  = ram_conduit_writedata[4];

assign \ram_conduit_writedata[5]~input_o  = ram_conduit_writedata[5];

assign \ram_conduit_writedata[6]~input_o  = ram_conduit_writedata[6];

assign \ram_conduit_writedata[7]~input_o  = ram_conduit_writedata[7];

assign \ram_conduit_writedata[8]~input_o  = ram_conduit_writedata[8];

assign \ram_conduit_byteenable[1]~input_o  = ram_conduit_byteenable[1];

assign \ram_conduit_writedata[9]~input_o  = ram_conduit_writedata[9];

assign \ram_conduit_writedata[10]~input_o  = ram_conduit_writedata[10];

assign \ram_conduit_writedata[11]~input_o  = ram_conduit_writedata[11];

assign \ram_conduit_writedata[12]~input_o  = ram_conduit_writedata[12];

assign \ram_conduit_writedata[13]~input_o  = ram_conduit_writedata[13];

assign \ram_conduit_writedata[14]~input_o  = ram_conduit_writedata[14];

assign \ram_conduit_writedata[15]~input_o  = ram_conduit_writedata[15];

assign \reset_reset_n~input_o  = reset_reset_n;

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck_n),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output (
	.i(\hps_0|hps_io|border|intermediate[36] ),
	.oe(\hps_0|hps_io|border|intermediate[37] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_spim1_inst_MOSI),
	.obar());
defparam \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .shift_series_termination_control = "false";

assign hps_io_hps_io_emac1_inst_TX_CLK = \hps_0|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;

assign hps_io_hps_io_emac1_inst_TXD0 = \hps_0|hps_io|border|emac1_inst~emac_phy_txd ;

assign hps_io_hps_io_emac1_inst_TXD1 = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;

assign hps_io_hps_io_emac1_inst_TXD2 = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;

assign hps_io_hps_io_emac1_inst_TXD3 = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;

assign hps_io_hps_io_emac1_inst_MDC = \hps_0|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;

assign hps_io_hps_io_emac1_inst_TX_CTL = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;

assign hps_io_hps_io_qspi_inst_SS0 = \hps_0|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;

assign hps_io_hps_io_qspi_inst_CLK = \hps_0|hps_io|border|qspi_inst~O_QSPI_SCLK ;

assign hps_io_hps_io_sdio_inst_CLK = \hps_0|hps_io|border|sdio_inst~sdmmc_cclk ;

assign hps_io_hps_io_usb1_inst_STP = \hps_0|hps_io|border|usb1_inst~usb_ulpi_stp ;

assign hps_io_hps_io_spim1_inst_CLK = \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;

assign hps_io_hps_io_spim1_inst_SS0 = \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;

assign hps_io_hps_io_uart0_inst_TX = \hps_0|hps_io|border|uart0_inst~uart_txd ;

assign memory_mem_a[0] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;

assign memory_mem_a[1] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;

assign memory_mem_a[2] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;

assign memory_mem_a[3] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;

assign memory_mem_a[4] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;

assign memory_mem_a[5] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;

assign memory_mem_a[6] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;

assign memory_mem_a[7] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;

assign memory_mem_a[8] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;

assign memory_mem_a[9] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;

assign memory_mem_a[10] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;

assign memory_mem_a[11] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;

assign memory_mem_a[12] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;

assign memory_mem_a[13] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;

assign memory_mem_a[14] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;

assign memory_mem_ba[0] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;

assign memory_mem_ba[1] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;

assign memory_mem_ba[2] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;

assign memory_mem_cke = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;

assign memory_mem_cs_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;

assign memory_mem_ras_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;

assign memory_mem_cas_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;

assign memory_mem_we_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;

assign memory_mem_reset_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;

assign memory_mem_odt = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;

assign ram_conduit_readdata[0] = \ram|the_altsyncram|auto_generated|q_b[0] ;

assign ram_conduit_readdata[1] = \ram|the_altsyncram|auto_generated|q_b[1] ;

assign ram_conduit_readdata[2] = \ram|the_altsyncram|auto_generated|q_b[2] ;

assign ram_conduit_readdata[3] = \ram|the_altsyncram|auto_generated|q_b[3] ;

assign ram_conduit_readdata[4] = \ram|the_altsyncram|auto_generated|q_b[4] ;

assign ram_conduit_readdata[5] = \ram|the_altsyncram|auto_generated|q_b[5] ;

assign ram_conduit_readdata[6] = \ram|the_altsyncram|auto_generated|q_b[6] ;

assign ram_conduit_readdata[7] = \ram|the_altsyncram|auto_generated|q_b[7] ;

assign ram_conduit_readdata[8] = \ram|the_altsyncram|auto_generated|q_b[8] ;

assign ram_conduit_readdata[9] = \ram|the_altsyncram|auto_generated|q_b[9] ;

assign ram_conduit_readdata[10] = \ram|the_altsyncram|auto_generated|q_b[10] ;

assign ram_conduit_readdata[11] = \ram|the_altsyncram|auto_generated|q_b[11] ;

assign ram_conduit_readdata[12] = \ram|the_altsyncram|auto_generated|q_b[12] ;

assign ram_conduit_readdata[13] = \ram|the_altsyncram|auto_generated|q_b[13] ;

assign ram_conduit_readdata[14] = \ram|the_altsyncram|auto_generated|q_b[14] ;

assign ram_conduit_readdata[15] = \ram|the_altsyncram|auto_generated|q_b[15] ;

assign vga_clk_ext_clk = \pll_0|altera_pll_i|outclk_wire[1] ;

assign vga_clk_int_clk = \pll_0|altera_pll_i|outclk_wire[0] ;

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output (
	.i(\hps_0|hps_io|border|intermediate[0] ),
	.oe(\hps_0|hps_io|border|intermediate[1] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_emac1_inst_MDIO),
	.obar());
defparam \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output (
	.i(\hps_0|hps_io|border|intermediate[2] ),
	.oe(\hps_0|hps_io|border|intermediate[3] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO0),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output (
	.i(\hps_0|hps_io|border|intermediate[4] ),
	.oe(\hps_0|hps_io|border|intermediate[5] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO1),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output (
	.i(\hps_0|hps_io|border|intermediate[6] ),
	.oe(\hps_0|hps_io|border|intermediate[7] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO2),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output (
	.i(\hps_0|hps_io|border|intermediate[8] ),
	.oe(\hps_0|hps_io|border|intermediate[9] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO3),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output (
	.i(\hps_0|hps_io|border|intermediate[10] ),
	.oe(\hps_0|hps_io|border|intermediate[11] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_CMD),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output (
	.i(\hps_0|hps_io|border|intermediate[12] ),
	.oe(\hps_0|hps_io|border|intermediate[13] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D0),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output (
	.i(\hps_0|hps_io|border|intermediate[14] ),
	.oe(\hps_0|hps_io|border|intermediate[15] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D1),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output (
	.i(\hps_0|hps_io|border|intermediate[16] ),
	.oe(\hps_0|hps_io|border|intermediate[17] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D2),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output (
	.i(\hps_0|hps_io|border|intermediate[18] ),
	.oe(\hps_0|hps_io|border|intermediate[19] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D3),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output (
	.i(\hps_0|hps_io|border|intermediate[20] ),
	.oe(\hps_0|hps_io|border|intermediate[21] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D0),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output (
	.i(\hps_0|hps_io|border|intermediate[22] ),
	.oe(\hps_0|hps_io|border|intermediate[23] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D1),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output (
	.i(\hps_0|hps_io|border|intermediate[24] ),
	.oe(\hps_0|hps_io|border|intermediate[25] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D2),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output (
	.i(\hps_0|hps_io|border|intermediate[26] ),
	.oe(\hps_0|hps_io|border|intermediate[27] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D3),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output (
	.i(\hps_0|hps_io|border|intermediate[28] ),
	.oe(\hps_0|hps_io|border|intermediate[29] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D4),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output (
	.i(\hps_0|hps_io|border|intermediate[30] ),
	.oe(\hps_0|hps_io|border|intermediate[31] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D5),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output (
	.i(\hps_0|hps_io|border|intermediate[32] ),
	.oe(\hps_0|hps_io|border|intermediate[33] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D6),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output (
	.i(\hps_0|hps_io|border|intermediate[34] ),
	.oe(\hps_0|hps_io|border|intermediate[35] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D7),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~output (
	.i(!\hps_0|hps_io|border|intermediate[38] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c0_inst_SDA),
	.obar());
defparam \hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .open_drain_output = "true";
defparam \hps_0|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~output (
	.i(!\hps_0|hps_io|border|intermediate[39] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c0_inst_SCL),
	.obar());
defparam \hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .open_drain_output = "true";
defparam \hps_0|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~output (
	.i(!\hps_0|hps_io|border|intermediate[40] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c1_inst_SDA),
	.obar());
defparam \hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .open_drain_output = "true";
defparam \hps_0|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~output (
	.i(!\hps_0|hps_io|border|intermediate[41] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c1_inst_SCL),
	.obar());
defparam \hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .open_drain_output = "true";
defparam \hps_0|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[4]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[5]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[6]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[7]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[8]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[9]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[10]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[11]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[12]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[13]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[14]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[15]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[16]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[17]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[18]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[19]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[20]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[21]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[22]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[23]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[24]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[25]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[26]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[27]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[28]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[29]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[30]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[31]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

endmodule

module system_altera_reset_controller (
	h2f_rst_n_0,
	merged_reset,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	merged_reset;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \merged_reset~0 (
	.dataa(!h2f_rst_n_0),
	.datab(!reset_reset_n),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(merged_reset),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_reset~0 .extended_lut = "off";
defparam \merged_reset~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \merged_reset~0 .shared_arith = "off";

endmodule

module system_altera_reset_controller_1 (
	r_early_rst1,
	merged_reset,
	r_sync_rst1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	r_early_rst1;
input 	merged_reset;
output 	r_sync_rst1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \always2~0_combout ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;


system_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk));

system_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.merged_reset(merged_reset),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk));

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h7373737373737373;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module system_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module system_altera_reset_synchronizer_1 (
	merged_reset,
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	merged_reset;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module system_altera_reset_controller_2 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.h2f_rst_n_0(h2f_rst_n_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

endmodule

module system_altera_reset_synchronizer_3 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module system_system_hps_0 (
	h2f_rst_n_0,
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	sink1_ready,
	awready,
	src0_valid,
	source_endofpacket,
	src1_valid,
	wready,
	mem_70_0,
	mem_71_0,
	mem_72_0,
	mem_73_0,
	mem_74_0,
	mem_75_0,
	mem_76_0,
	mem_77_0,
	mem_78_0,
	mem_79_0,
	mem_80_0,
	mem_81_0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	ShiftLeft2,
	ShiftLeft21,
	ShiftLeft22,
	ShiftLeft23,
	ShiftLeft24,
	ShiftLeft25,
	ShiftLeft26,
	ShiftLeft27,
	ShiftLeft28,
	ShiftLeft29,
	ShiftLeft210,
	ShiftLeft211,
	ShiftLeft212,
	ShiftLeft213,
	ShiftLeft214,
	ShiftLeft215,
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim1_inst,
	spim1_inst1,
	intermediate_36,
	intermediate_37,
	uart0_inst,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	clk_clk,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	h2f_rst_n_0;
output 	h2f_lw_ARVALID_0;
output 	h2f_lw_AWVALID_0;
output 	h2f_lw_BREADY_0;
output 	h2f_lw_RREADY_0;
output 	h2f_lw_WLAST_0;
output 	h2f_lw_WVALID_0;
output 	h2f_lw_ARADDR_0;
output 	h2f_lw_ARADDR_1;
output 	h2f_lw_ARADDR_2;
output 	h2f_lw_ARADDR_3;
output 	h2f_lw_ARADDR_4;
output 	h2f_lw_ARBURST_0;
output 	h2f_lw_ARBURST_1;
output 	h2f_lw_ARID_0;
output 	h2f_lw_ARID_1;
output 	h2f_lw_ARID_2;
output 	h2f_lw_ARID_3;
output 	h2f_lw_ARID_4;
output 	h2f_lw_ARID_5;
output 	h2f_lw_ARID_6;
output 	h2f_lw_ARID_7;
output 	h2f_lw_ARID_8;
output 	h2f_lw_ARID_9;
output 	h2f_lw_ARID_10;
output 	h2f_lw_ARID_11;
output 	h2f_lw_ARLEN_0;
output 	h2f_lw_ARLEN_1;
output 	h2f_lw_ARLEN_2;
output 	h2f_lw_ARLEN_3;
output 	h2f_lw_ARSIZE_0;
output 	h2f_lw_ARSIZE_1;
output 	h2f_lw_ARSIZE_2;
output 	h2f_lw_AWADDR_0;
output 	h2f_lw_AWADDR_1;
output 	h2f_lw_AWADDR_2;
output 	h2f_lw_AWADDR_3;
output 	h2f_lw_AWADDR_4;
output 	h2f_lw_AWBURST_0;
output 	h2f_lw_AWBURST_1;
output 	h2f_lw_AWID_0;
output 	h2f_lw_AWID_1;
output 	h2f_lw_AWID_2;
output 	h2f_lw_AWID_3;
output 	h2f_lw_AWID_4;
output 	h2f_lw_AWID_5;
output 	h2f_lw_AWID_6;
output 	h2f_lw_AWID_7;
output 	h2f_lw_AWID_8;
output 	h2f_lw_AWID_9;
output 	h2f_lw_AWID_10;
output 	h2f_lw_AWID_11;
output 	h2f_lw_AWLEN_0;
output 	h2f_lw_AWLEN_1;
output 	h2f_lw_AWLEN_2;
output 	h2f_lw_AWLEN_3;
output 	h2f_lw_AWSIZE_0;
output 	h2f_lw_AWSIZE_1;
output 	h2f_lw_AWSIZE_2;
output 	h2f_lw_WDATA_0;
output 	h2f_lw_WDATA_1;
output 	h2f_lw_WDATA_2;
output 	h2f_lw_WDATA_3;
output 	h2f_lw_WDATA_4;
output 	h2f_lw_WDATA_5;
output 	h2f_lw_WDATA_6;
output 	h2f_lw_WDATA_7;
output 	h2f_lw_WDATA_8;
output 	h2f_lw_WDATA_9;
output 	h2f_lw_WDATA_10;
output 	h2f_lw_WDATA_11;
output 	h2f_lw_WDATA_12;
output 	h2f_lw_WDATA_13;
output 	h2f_lw_WDATA_14;
output 	h2f_lw_WDATA_15;
output 	h2f_lw_WDATA_16;
output 	h2f_lw_WDATA_17;
output 	h2f_lw_WDATA_18;
output 	h2f_lw_WDATA_19;
output 	h2f_lw_WDATA_20;
output 	h2f_lw_WDATA_21;
output 	h2f_lw_WDATA_22;
output 	h2f_lw_WDATA_23;
output 	h2f_lw_WDATA_24;
output 	h2f_lw_WDATA_25;
output 	h2f_lw_WDATA_26;
output 	h2f_lw_WDATA_27;
output 	h2f_lw_WDATA_28;
output 	h2f_lw_WDATA_29;
output 	h2f_lw_WDATA_30;
output 	h2f_lw_WDATA_31;
output 	h2f_lw_WSTRB_0;
output 	h2f_lw_WSTRB_1;
output 	h2f_lw_WSTRB_2;
output 	h2f_lw_WSTRB_3;
input 	sink1_ready;
input 	awready;
input 	src0_valid;
input 	source_endofpacket;
input 	src1_valid;
input 	wready;
input 	mem_70_0;
input 	mem_71_0;
input 	mem_72_0;
input 	mem_73_0;
input 	mem_74_0;
input 	mem_75_0;
input 	mem_76_0;
input 	mem_77_0;
input 	mem_78_0;
input 	mem_79_0;
input 	mem_80_0;
input 	mem_81_0;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	out_data_8;
input 	out_data_9;
input 	out_data_10;
input 	out_data_11;
input 	out_data_12;
input 	out_data_13;
input 	out_data_14;
input 	out_data_15;
input 	ShiftLeft2;
input 	ShiftLeft21;
input 	ShiftLeft22;
input 	ShiftLeft23;
input 	ShiftLeft24;
input 	ShiftLeft25;
input 	ShiftLeft26;
input 	ShiftLeft27;
input 	ShiftLeft28;
input 	ShiftLeft29;
input 	ShiftLeft210;
input 	ShiftLeft211;
input 	ShiftLeft212;
input 	ShiftLeft213;
input 	ShiftLeft214;
input 	ShiftLeft215;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	uart0_inst;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	clk_clk;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_system_hps_0_hps_io hps_io(
	.emac1_inst(emac1_inst),
	.emac1_inst1(emac1_inst1),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.emac1_inst2(emac1_inst2),
	.emac1_inst3(emac1_inst3),
	.emac1_inst4(emac1_inst4),
	.emac1_inst5(emac1_inst5),
	.emac1_inst6(emac1_inst6),
	.qspi_inst(qspi_inst),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.qspi_inst1(qspi_inst1),
	.sdio_inst(sdio_inst),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.usb1_inst(usb1_inst),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.spim1_inst(spim1_inst),
	.spim1_inst1(spim1_inst1),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.uart0_inst(uart0_inst),
	.intermediate_39(intermediate_39),
	.intermediate_38(intermediate_38),
	.intermediate_41(intermediate_41),
	.intermediate_40(intermediate_40),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_i2c0_inst_SDA_0(hps_io_i2c0_inst_SDA_0),
	.hps_io_i2c0_inst_SCL_0(hps_io_i2c0_inst_SCL_0),
	.hps_io_i2c1_inst_SDA_0(hps_io_i2c1_inst_SDA_0),
	.hps_io_i2c1_inst_SCL_0(hps_io_i2c1_inst_SCL_0),
	.hps_io_hps_io_emac1_inst_RXD0(hps_io_hps_io_emac1_inst_RXD0),
	.hps_io_hps_io_emac1_inst_RXD1(hps_io_hps_io_emac1_inst_RXD1),
	.hps_io_hps_io_emac1_inst_RXD2(hps_io_hps_io_emac1_inst_RXD2),
	.hps_io_hps_io_emac1_inst_RXD3(hps_io_hps_io_emac1_inst_RXD3),
	.hps_io_hps_io_emac1_inst_RX_CLK(hps_io_hps_io_emac1_inst_RX_CLK),
	.hps_io_hps_io_emac1_inst_RX_CTL(hps_io_hps_io_emac1_inst_RX_CTL),
	.hps_io_hps_io_spim1_inst_MISO(hps_io_hps_io_spim1_inst_MISO),
	.hps_io_hps_io_uart0_inst_RX(hps_io_hps_io_uart0_inst_RX),
	.hps_io_hps_io_usb1_inst_CLK(hps_io_hps_io_usb1_inst_CLK),
	.hps_io_hps_io_usb1_inst_DIR(hps_io_hps_io_usb1_inst_DIR),
	.hps_io_hps_io_usb1_inst_NXT(hps_io_hps_io_usb1_inst_NXT),
	.memory_oct_rzqin(memory_oct_rzqin));

system_system_hps_0_fpga_interfaces fpga_interfaces(
	.h2f_rst_n({h2f_rst_n_0}),
	.h2f_lw_ARVALID({h2f_lw_ARVALID_0}),
	.h2f_lw_AWVALID({h2f_lw_AWVALID_0}),
	.h2f_lw_BREADY({h2f_lw_BREADY_0}),
	.h2f_lw_RREADY({h2f_lw_RREADY_0}),
	.h2f_lw_WLAST({h2f_lw_WLAST_0}),
	.h2f_lw_WVALID({h2f_lw_WVALID_0}),
	.h2f_lw_ARADDR({h2f_lw_ARADDR_unconnected_wire_20,h2f_lw_ARADDR_unconnected_wire_19,h2f_lw_ARADDR_unconnected_wire_18,h2f_lw_ARADDR_unconnected_wire_17,h2f_lw_ARADDR_unconnected_wire_16,h2f_lw_ARADDR_unconnected_wire_15,h2f_lw_ARADDR_unconnected_wire_14,
h2f_lw_ARADDR_unconnected_wire_13,h2f_lw_ARADDR_unconnected_wire_12,h2f_lw_ARADDR_unconnected_wire_11,h2f_lw_ARADDR_unconnected_wire_10,h2f_lw_ARADDR_unconnected_wire_9,h2f_lw_ARADDR_unconnected_wire_8,h2f_lw_ARADDR_unconnected_wire_7,
h2f_lw_ARADDR_unconnected_wire_6,h2f_lw_ARADDR_unconnected_wire_5,h2f_lw_ARADDR_4,h2f_lw_ARADDR_3,h2f_lw_ARADDR_2,h2f_lw_ARADDR_1,h2f_lw_ARADDR_0}),
	.h2f_lw_ARBURST({h2f_lw_ARBURST_1,h2f_lw_ARBURST_0}),
	.h2f_lw_ARID({h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0}),
	.h2f_lw_ARLEN({h2f_lw_ARLEN_3,h2f_lw_ARLEN_2,h2f_lw_ARLEN_1,h2f_lw_ARLEN_0}),
	.h2f_lw_ARSIZE({h2f_lw_ARSIZE_2,h2f_lw_ARSIZE_1,h2f_lw_ARSIZE_0}),
	.h2f_lw_AWADDR({h2f_lw_AWADDR_unconnected_wire_20,h2f_lw_AWADDR_unconnected_wire_19,h2f_lw_AWADDR_unconnected_wire_18,h2f_lw_AWADDR_unconnected_wire_17,h2f_lw_AWADDR_unconnected_wire_16,h2f_lw_AWADDR_unconnected_wire_15,h2f_lw_AWADDR_unconnected_wire_14,
h2f_lw_AWADDR_unconnected_wire_13,h2f_lw_AWADDR_unconnected_wire_12,h2f_lw_AWADDR_unconnected_wire_11,h2f_lw_AWADDR_unconnected_wire_10,h2f_lw_AWADDR_unconnected_wire_9,h2f_lw_AWADDR_unconnected_wire_8,h2f_lw_AWADDR_unconnected_wire_7,
h2f_lw_AWADDR_unconnected_wire_6,h2f_lw_AWADDR_unconnected_wire_5,h2f_lw_AWADDR_4,h2f_lw_AWADDR_3,h2f_lw_AWADDR_2,h2f_lw_AWADDR_1,h2f_lw_AWADDR_0}),
	.h2f_lw_AWBURST({h2f_lw_AWBURST_1,h2f_lw_AWBURST_0}),
	.h2f_lw_AWID({h2f_lw_AWID_11,h2f_lw_AWID_10,h2f_lw_AWID_9,h2f_lw_AWID_8,h2f_lw_AWID_7,h2f_lw_AWID_6,h2f_lw_AWID_5,h2f_lw_AWID_4,h2f_lw_AWID_3,h2f_lw_AWID_2,h2f_lw_AWID_1,h2f_lw_AWID_0}),
	.h2f_lw_AWLEN({h2f_lw_AWLEN_3,h2f_lw_AWLEN_2,h2f_lw_AWLEN_1,h2f_lw_AWLEN_0}),
	.h2f_lw_AWSIZE({h2f_lw_AWSIZE_2,h2f_lw_AWSIZE_1,h2f_lw_AWSIZE_0}),
	.h2f_lw_WDATA({h2f_lw_WDATA_31,h2f_lw_WDATA_30,h2f_lw_WDATA_29,h2f_lw_WDATA_28,h2f_lw_WDATA_27,h2f_lw_WDATA_26,h2f_lw_WDATA_25,h2f_lw_WDATA_24,h2f_lw_WDATA_23,h2f_lw_WDATA_22,h2f_lw_WDATA_21,h2f_lw_WDATA_20,h2f_lw_WDATA_19,h2f_lw_WDATA_18,h2f_lw_WDATA_17,h2f_lw_WDATA_16,h2f_lw_WDATA_15,
h2f_lw_WDATA_14,h2f_lw_WDATA_13,h2f_lw_WDATA_12,h2f_lw_WDATA_11,h2f_lw_WDATA_10,h2f_lw_WDATA_9,h2f_lw_WDATA_8,h2f_lw_WDATA_7,h2f_lw_WDATA_6,h2f_lw_WDATA_5,h2f_lw_WDATA_4,h2f_lw_WDATA_3,h2f_lw_WDATA_2,h2f_lw_WDATA_1,h2f_lw_WDATA_0}),
	.h2f_lw_WSTRB({h2f_lw_WSTRB_3,h2f_lw_WSTRB_2,h2f_lw_WSTRB_1,h2f_lw_WSTRB_0}),
	.h2f_lw_ARREADY({sink1_ready}),
	.h2f_lw_AWREADY({awready}),
	.h2f_lw_BVALID({src0_valid}),
	.h2f_lw_RLAST({source_endofpacket}),
	.h2f_lw_RVALID({src1_valid}),
	.h2f_lw_WREADY({wready}),
	.h2f_lw_BID({mem_81_0,mem_80_0,mem_79_0,mem_78_0,mem_77_0,mem_76_0,mem_75_0,mem_74_0,mem_73_0,mem_72_0,mem_71_0,mem_70_0}),
	.h2f_lw_RID({mem_81_0,mem_80_0,mem_79_0,mem_78_0,mem_77_0,mem_76_0,mem_75_0,mem_74_0,mem_73_0,mem_72_0,mem_71_0,mem_70_0}),
	.h2f_lw_RDATA({ShiftLeft215,ShiftLeft214,ShiftLeft213,ShiftLeft212,ShiftLeft211,ShiftLeft210,ShiftLeft29,ShiftLeft28,ShiftLeft27,ShiftLeft26,ShiftLeft25,ShiftLeft24,ShiftLeft23,ShiftLeft22,ShiftLeft21,ShiftLeft2,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,out_data_10,
out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.f2h_axi_clk({clk_clk}),
	.h2f_axi_clk({clk_clk}),
	.h2f_lw_axi_clk({clk_clk}));

endmodule

module system_system_hps_0_fpga_interfaces (
	h2f_rst_n,
	h2f_lw_ARVALID,
	h2f_lw_AWVALID,
	h2f_lw_BREADY,
	h2f_lw_RREADY,
	h2f_lw_WLAST,
	h2f_lw_WVALID,
	h2f_lw_ARADDR,
	h2f_lw_ARBURST,
	h2f_lw_ARID,
	h2f_lw_ARLEN,
	h2f_lw_ARSIZE,
	h2f_lw_AWADDR,
	h2f_lw_AWBURST,
	h2f_lw_AWID,
	h2f_lw_AWLEN,
	h2f_lw_AWSIZE,
	h2f_lw_WDATA,
	h2f_lw_WSTRB,
	h2f_lw_ARREADY,
	h2f_lw_AWREADY,
	h2f_lw_BVALID,
	h2f_lw_RLAST,
	h2f_lw_RVALID,
	h2f_lw_WREADY,
	h2f_lw_BID,
	h2f_lw_RID,
	h2f_lw_RDATA,
	f2h_axi_clk,
	h2f_axi_clk,
	h2f_lw_axi_clk)/* synthesis synthesis_greybox=0 */;
output 	[0:0] h2f_rst_n;
output 	[0:0] h2f_lw_ARVALID;
output 	[0:0] h2f_lw_AWVALID;
output 	[0:0] h2f_lw_BREADY;
output 	[0:0] h2f_lw_RREADY;
output 	[0:0] h2f_lw_WLAST;
output 	[0:0] h2f_lw_WVALID;
output 	[20:0] h2f_lw_ARADDR;
output 	[1:0] h2f_lw_ARBURST;
output 	[11:0] h2f_lw_ARID;
output 	[3:0] h2f_lw_ARLEN;
output 	[2:0] h2f_lw_ARSIZE;
output 	[20:0] h2f_lw_AWADDR;
output 	[1:0] h2f_lw_AWBURST;
output 	[11:0] h2f_lw_AWID;
output 	[3:0] h2f_lw_AWLEN;
output 	[2:0] h2f_lw_AWSIZE;
output 	[31:0] h2f_lw_WDATA;
output 	[3:0] h2f_lw_WSTRB;
input 	[0:0] h2f_lw_ARREADY;
input 	[0:0] h2f_lw_AWREADY;
input 	[0:0] h2f_lw_BVALID;
input 	[0:0] h2f_lw_RLAST;
input 	[0:0] h2f_lw_RVALID;
input 	[0:0] h2f_lw_WREADY;
input 	[11:0] h2f_lw_BID;
input 	[11:0] h2f_lw_RID;
input 	[31:0] h2f_lw_RDATA;
input 	[0:0] f2h_axi_clk;
input 	[0:0] h2f_axi_clk;
input 	[0:0] h2f_lw_axi_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \debug_apb~O_P_ADDR_31 ;
wire \tpiu~trace_data ;
wire \tpiu~O_TRACE_DATA1 ;
wire \tpiu~O_TRACE_DATA2 ;
wire \tpiu~O_TRACE_DATA3 ;
wire \tpiu~O_TRACE_DATA4 ;
wire \tpiu~O_TRACE_DATA5 ;
wire \tpiu~O_TRACE_DATA6 ;
wire \tpiu~O_TRACE_DATA7 ;
wire \tpiu~O_TRACE_DATA8 ;
wire \tpiu~O_TRACE_DATA9 ;
wire \tpiu~O_TRACE_DATA10 ;
wire \tpiu~O_TRACE_DATA11 ;
wire \tpiu~O_TRACE_DATA12 ;
wire \tpiu~O_TRACE_DATA13 ;
wire \tpiu~O_TRACE_DATA14 ;
wire \tpiu~O_TRACE_DATA15 ;
wire \tpiu~O_TRACE_DATA16 ;
wire \tpiu~O_TRACE_DATA17 ;
wire \tpiu~O_TRACE_DATA18 ;
wire \tpiu~O_TRACE_DATA19 ;
wire \tpiu~O_TRACE_DATA20 ;
wire \tpiu~O_TRACE_DATA21 ;
wire \tpiu~O_TRACE_DATA22 ;
wire \tpiu~O_TRACE_DATA23 ;
wire \tpiu~O_TRACE_DATA24 ;
wire \tpiu~O_TRACE_DATA25 ;
wire \tpiu~O_TRACE_DATA26 ;
wire \tpiu~O_TRACE_DATA27 ;
wire \tpiu~O_TRACE_DATA28 ;
wire \tpiu~O_TRACE_DATA29 ;
wire \tpiu~O_TRACE_DATA30 ;
wire \tpiu~O_TRACE_DATA31 ;
wire \boot_from_fpga~fake_dout ;
wire \f2h_ARREADY[0] ;
wire \h2f_ARADDR[0] ;
wire \h2f_ARADDR[1] ;
wire \h2f_ARADDR[2] ;
wire \h2f_ARADDR[3] ;
wire \h2f_ARADDR[4] ;
wire \h2f_ARADDR[5] ;
wire \h2f_ARADDR[6] ;
wire \h2f_ARADDR[7] ;
wire \h2f_ARADDR[8] ;
wire \h2f_ARADDR[9] ;
wire \h2f_ARADDR[10] ;
wire \h2f_ARADDR[11] ;
wire \h2f_ARADDR[12] ;
wire \h2f_ARADDR[13] ;
wire \h2f_ARADDR[14] ;
wire \h2f_ARADDR[15] ;
wire \h2f_ARADDR[16] ;
wire \h2f_ARADDR[17] ;
wire \h2f_ARADDR[18] ;
wire \h2f_ARADDR[19] ;
wire \h2f_ARADDR[20] ;
wire \h2f_ARADDR[21] ;
wire \h2f_ARADDR[22] ;
wire \h2f_ARADDR[23] ;
wire \h2f_ARADDR[24] ;
wire \h2f_ARADDR[25] ;
wire \h2f_ARADDR[26] ;
wire \h2f_ARADDR[27] ;
wire \h2f_ARADDR[28] ;
wire \h2f_ARADDR[29] ;
wire \f2sdram~O_BONDING_OUT_10 ;
wire \f2sdram~O_BONDING_OUT_11 ;
wire \f2sdram~O_BONDING_OUT_12 ;
wire \f2sdram~O_BONDING_OUT_13 ;
wire \interrupts~fake_dout ;
wire \clocks_resets~h2f_cold_rst_n ;
wire \h2f_lw_ARADDR[5] ;
wire \h2f_lw_ARADDR[6] ;
wire \h2f_lw_ARADDR[7] ;
wire \h2f_lw_ARADDR[8] ;
wire \h2f_lw_ARADDR[9] ;
wire \h2f_lw_ARADDR[10] ;
wire \h2f_lw_ARADDR[11] ;
wire \h2f_lw_ARADDR[12] ;
wire \h2f_lw_ARADDR[13] ;
wire \h2f_lw_ARADDR[14] ;
wire \h2f_lw_ARADDR[15] ;
wire \h2f_lw_ARADDR[16] ;
wire \h2f_lw_ARADDR[17] ;
wire \h2f_lw_ARADDR[18] ;
wire \h2f_lw_ARADDR[19] ;
wire \h2f_lw_ARADDR[20] ;

wire [31:0] tpiu_TRACE_DATA_bus;
wire [29:0] hps2fpga_ARADDR_bus;
wire [3:0] f2sdram_BONDING_OUT_1_bus;
wire [20:0] hps2fpga_light_weight_ARADDR_bus;
wire [1:0] hps2fpga_light_weight_ARBURST_bus;
wire [11:0] hps2fpga_light_weight_ARID_bus;
wire [3:0] hps2fpga_light_weight_ARLEN_bus;
wire [2:0] hps2fpga_light_weight_ARSIZE_bus;
wire [20:0] hps2fpga_light_weight_AWADDR_bus;
wire [1:0] hps2fpga_light_weight_AWBURST_bus;
wire [11:0] hps2fpga_light_weight_AWID_bus;
wire [3:0] hps2fpga_light_weight_AWLEN_bus;
wire [2:0] hps2fpga_light_weight_AWSIZE_bus;
wire [31:0] hps2fpga_light_weight_WDATA_bus;
wire [3:0] hps2fpga_light_weight_WSTRB_bus;

assign \tpiu~trace_data  = tpiu_TRACE_DATA_bus[0];
assign \tpiu~O_TRACE_DATA1  = tpiu_TRACE_DATA_bus[1];
assign \tpiu~O_TRACE_DATA2  = tpiu_TRACE_DATA_bus[2];
assign \tpiu~O_TRACE_DATA3  = tpiu_TRACE_DATA_bus[3];
assign \tpiu~O_TRACE_DATA4  = tpiu_TRACE_DATA_bus[4];
assign \tpiu~O_TRACE_DATA5  = tpiu_TRACE_DATA_bus[5];
assign \tpiu~O_TRACE_DATA6  = tpiu_TRACE_DATA_bus[6];
assign \tpiu~O_TRACE_DATA7  = tpiu_TRACE_DATA_bus[7];
assign \tpiu~O_TRACE_DATA8  = tpiu_TRACE_DATA_bus[8];
assign \tpiu~O_TRACE_DATA9  = tpiu_TRACE_DATA_bus[9];
assign \tpiu~O_TRACE_DATA10  = tpiu_TRACE_DATA_bus[10];
assign \tpiu~O_TRACE_DATA11  = tpiu_TRACE_DATA_bus[11];
assign \tpiu~O_TRACE_DATA12  = tpiu_TRACE_DATA_bus[12];
assign \tpiu~O_TRACE_DATA13  = tpiu_TRACE_DATA_bus[13];
assign \tpiu~O_TRACE_DATA14  = tpiu_TRACE_DATA_bus[14];
assign \tpiu~O_TRACE_DATA15  = tpiu_TRACE_DATA_bus[15];
assign \tpiu~O_TRACE_DATA16  = tpiu_TRACE_DATA_bus[16];
assign \tpiu~O_TRACE_DATA17  = tpiu_TRACE_DATA_bus[17];
assign \tpiu~O_TRACE_DATA18  = tpiu_TRACE_DATA_bus[18];
assign \tpiu~O_TRACE_DATA19  = tpiu_TRACE_DATA_bus[19];
assign \tpiu~O_TRACE_DATA20  = tpiu_TRACE_DATA_bus[20];
assign \tpiu~O_TRACE_DATA21  = tpiu_TRACE_DATA_bus[21];
assign \tpiu~O_TRACE_DATA22  = tpiu_TRACE_DATA_bus[22];
assign \tpiu~O_TRACE_DATA23  = tpiu_TRACE_DATA_bus[23];
assign \tpiu~O_TRACE_DATA24  = tpiu_TRACE_DATA_bus[24];
assign \tpiu~O_TRACE_DATA25  = tpiu_TRACE_DATA_bus[25];
assign \tpiu~O_TRACE_DATA26  = tpiu_TRACE_DATA_bus[26];
assign \tpiu~O_TRACE_DATA27  = tpiu_TRACE_DATA_bus[27];
assign \tpiu~O_TRACE_DATA28  = tpiu_TRACE_DATA_bus[28];
assign \tpiu~O_TRACE_DATA29  = tpiu_TRACE_DATA_bus[29];
assign \tpiu~O_TRACE_DATA30  = tpiu_TRACE_DATA_bus[30];
assign \tpiu~O_TRACE_DATA31  = tpiu_TRACE_DATA_bus[31];

assign \h2f_ARADDR[0]  = hps2fpga_ARADDR_bus[0];
assign \h2f_ARADDR[1]  = hps2fpga_ARADDR_bus[1];
assign \h2f_ARADDR[2]  = hps2fpga_ARADDR_bus[2];
assign \h2f_ARADDR[3]  = hps2fpga_ARADDR_bus[3];
assign \h2f_ARADDR[4]  = hps2fpga_ARADDR_bus[4];
assign \h2f_ARADDR[5]  = hps2fpga_ARADDR_bus[5];
assign \h2f_ARADDR[6]  = hps2fpga_ARADDR_bus[6];
assign \h2f_ARADDR[7]  = hps2fpga_ARADDR_bus[7];
assign \h2f_ARADDR[8]  = hps2fpga_ARADDR_bus[8];
assign \h2f_ARADDR[9]  = hps2fpga_ARADDR_bus[9];
assign \h2f_ARADDR[10]  = hps2fpga_ARADDR_bus[10];
assign \h2f_ARADDR[11]  = hps2fpga_ARADDR_bus[11];
assign \h2f_ARADDR[12]  = hps2fpga_ARADDR_bus[12];
assign \h2f_ARADDR[13]  = hps2fpga_ARADDR_bus[13];
assign \h2f_ARADDR[14]  = hps2fpga_ARADDR_bus[14];
assign \h2f_ARADDR[15]  = hps2fpga_ARADDR_bus[15];
assign \h2f_ARADDR[16]  = hps2fpga_ARADDR_bus[16];
assign \h2f_ARADDR[17]  = hps2fpga_ARADDR_bus[17];
assign \h2f_ARADDR[18]  = hps2fpga_ARADDR_bus[18];
assign \h2f_ARADDR[19]  = hps2fpga_ARADDR_bus[19];
assign \h2f_ARADDR[20]  = hps2fpga_ARADDR_bus[20];
assign \h2f_ARADDR[21]  = hps2fpga_ARADDR_bus[21];
assign \h2f_ARADDR[22]  = hps2fpga_ARADDR_bus[22];
assign \h2f_ARADDR[23]  = hps2fpga_ARADDR_bus[23];
assign \h2f_ARADDR[24]  = hps2fpga_ARADDR_bus[24];
assign \h2f_ARADDR[25]  = hps2fpga_ARADDR_bus[25];
assign \h2f_ARADDR[26]  = hps2fpga_ARADDR_bus[26];
assign \h2f_ARADDR[27]  = hps2fpga_ARADDR_bus[27];
assign \h2f_ARADDR[28]  = hps2fpga_ARADDR_bus[28];
assign \h2f_ARADDR[29]  = hps2fpga_ARADDR_bus[29];

assign \f2sdram~O_BONDING_OUT_10  = f2sdram_BONDING_OUT_1_bus[0];
assign \f2sdram~O_BONDING_OUT_11  = f2sdram_BONDING_OUT_1_bus[1];
assign \f2sdram~O_BONDING_OUT_12  = f2sdram_BONDING_OUT_1_bus[2];
assign \f2sdram~O_BONDING_OUT_13  = f2sdram_BONDING_OUT_1_bus[3];

assign h2f_lw_ARADDR[0] = hps2fpga_light_weight_ARADDR_bus[0];
assign h2f_lw_ARADDR[1] = hps2fpga_light_weight_ARADDR_bus[1];
assign h2f_lw_ARADDR[2] = hps2fpga_light_weight_ARADDR_bus[2];
assign h2f_lw_ARADDR[3] = hps2fpga_light_weight_ARADDR_bus[3];
assign h2f_lw_ARADDR[4] = hps2fpga_light_weight_ARADDR_bus[4];
assign \h2f_lw_ARADDR[5]  = hps2fpga_light_weight_ARADDR_bus[5];
assign \h2f_lw_ARADDR[6]  = hps2fpga_light_weight_ARADDR_bus[6];
assign \h2f_lw_ARADDR[7]  = hps2fpga_light_weight_ARADDR_bus[7];
assign \h2f_lw_ARADDR[8]  = hps2fpga_light_weight_ARADDR_bus[8];
assign \h2f_lw_ARADDR[9]  = hps2fpga_light_weight_ARADDR_bus[9];
assign \h2f_lw_ARADDR[10]  = hps2fpga_light_weight_ARADDR_bus[10];
assign \h2f_lw_ARADDR[11]  = hps2fpga_light_weight_ARADDR_bus[11];
assign \h2f_lw_ARADDR[12]  = hps2fpga_light_weight_ARADDR_bus[12];
assign \h2f_lw_ARADDR[13]  = hps2fpga_light_weight_ARADDR_bus[13];
assign \h2f_lw_ARADDR[14]  = hps2fpga_light_weight_ARADDR_bus[14];
assign \h2f_lw_ARADDR[15]  = hps2fpga_light_weight_ARADDR_bus[15];
assign \h2f_lw_ARADDR[16]  = hps2fpga_light_weight_ARADDR_bus[16];
assign \h2f_lw_ARADDR[17]  = hps2fpga_light_weight_ARADDR_bus[17];
assign \h2f_lw_ARADDR[18]  = hps2fpga_light_weight_ARADDR_bus[18];
assign \h2f_lw_ARADDR[19]  = hps2fpga_light_weight_ARADDR_bus[19];
assign \h2f_lw_ARADDR[20]  = hps2fpga_light_weight_ARADDR_bus[20];

assign h2f_lw_ARBURST[0] = hps2fpga_light_weight_ARBURST_bus[0];
assign h2f_lw_ARBURST[1] = hps2fpga_light_weight_ARBURST_bus[1];

assign h2f_lw_ARID[0] = hps2fpga_light_weight_ARID_bus[0];
assign h2f_lw_ARID[1] = hps2fpga_light_weight_ARID_bus[1];
assign h2f_lw_ARID[2] = hps2fpga_light_weight_ARID_bus[2];
assign h2f_lw_ARID[3] = hps2fpga_light_weight_ARID_bus[3];
assign h2f_lw_ARID[4] = hps2fpga_light_weight_ARID_bus[4];
assign h2f_lw_ARID[5] = hps2fpga_light_weight_ARID_bus[5];
assign h2f_lw_ARID[6] = hps2fpga_light_weight_ARID_bus[6];
assign h2f_lw_ARID[7] = hps2fpga_light_weight_ARID_bus[7];
assign h2f_lw_ARID[8] = hps2fpga_light_weight_ARID_bus[8];
assign h2f_lw_ARID[9] = hps2fpga_light_weight_ARID_bus[9];
assign h2f_lw_ARID[10] = hps2fpga_light_weight_ARID_bus[10];
assign h2f_lw_ARID[11] = hps2fpga_light_weight_ARID_bus[11];

assign h2f_lw_ARLEN[0] = hps2fpga_light_weight_ARLEN_bus[0];
assign h2f_lw_ARLEN[1] = hps2fpga_light_weight_ARLEN_bus[1];
assign h2f_lw_ARLEN[2] = hps2fpga_light_weight_ARLEN_bus[2];
assign h2f_lw_ARLEN[3] = hps2fpga_light_weight_ARLEN_bus[3];

assign h2f_lw_ARSIZE[0] = hps2fpga_light_weight_ARSIZE_bus[0];
assign h2f_lw_ARSIZE[1] = hps2fpga_light_weight_ARSIZE_bus[1];
assign h2f_lw_ARSIZE[2] = hps2fpga_light_weight_ARSIZE_bus[2];

assign h2f_lw_AWADDR[0] = hps2fpga_light_weight_AWADDR_bus[0];
assign h2f_lw_AWADDR[1] = hps2fpga_light_weight_AWADDR_bus[1];
assign h2f_lw_AWADDR[2] = hps2fpga_light_weight_AWADDR_bus[2];
assign h2f_lw_AWADDR[3] = hps2fpga_light_weight_AWADDR_bus[3];
assign h2f_lw_AWADDR[4] = hps2fpga_light_weight_AWADDR_bus[4];

assign h2f_lw_AWBURST[0] = hps2fpga_light_weight_AWBURST_bus[0];
assign h2f_lw_AWBURST[1] = hps2fpga_light_weight_AWBURST_bus[1];

assign h2f_lw_AWID[0] = hps2fpga_light_weight_AWID_bus[0];
assign h2f_lw_AWID[1] = hps2fpga_light_weight_AWID_bus[1];
assign h2f_lw_AWID[2] = hps2fpga_light_weight_AWID_bus[2];
assign h2f_lw_AWID[3] = hps2fpga_light_weight_AWID_bus[3];
assign h2f_lw_AWID[4] = hps2fpga_light_weight_AWID_bus[4];
assign h2f_lw_AWID[5] = hps2fpga_light_weight_AWID_bus[5];
assign h2f_lw_AWID[6] = hps2fpga_light_weight_AWID_bus[6];
assign h2f_lw_AWID[7] = hps2fpga_light_weight_AWID_bus[7];
assign h2f_lw_AWID[8] = hps2fpga_light_weight_AWID_bus[8];
assign h2f_lw_AWID[9] = hps2fpga_light_weight_AWID_bus[9];
assign h2f_lw_AWID[10] = hps2fpga_light_weight_AWID_bus[10];
assign h2f_lw_AWID[11] = hps2fpga_light_weight_AWID_bus[11];

assign h2f_lw_AWLEN[0] = hps2fpga_light_weight_AWLEN_bus[0];
assign h2f_lw_AWLEN[1] = hps2fpga_light_weight_AWLEN_bus[1];
assign h2f_lw_AWLEN[2] = hps2fpga_light_weight_AWLEN_bus[2];
assign h2f_lw_AWLEN[3] = hps2fpga_light_weight_AWLEN_bus[3];

assign h2f_lw_AWSIZE[0] = hps2fpga_light_weight_AWSIZE_bus[0];
assign h2f_lw_AWSIZE[1] = hps2fpga_light_weight_AWSIZE_bus[1];
assign h2f_lw_AWSIZE[2] = hps2fpga_light_weight_AWSIZE_bus[2];

assign h2f_lw_WDATA[0] = hps2fpga_light_weight_WDATA_bus[0];
assign h2f_lw_WDATA[1] = hps2fpga_light_weight_WDATA_bus[1];
assign h2f_lw_WDATA[2] = hps2fpga_light_weight_WDATA_bus[2];
assign h2f_lw_WDATA[3] = hps2fpga_light_weight_WDATA_bus[3];
assign h2f_lw_WDATA[4] = hps2fpga_light_weight_WDATA_bus[4];
assign h2f_lw_WDATA[5] = hps2fpga_light_weight_WDATA_bus[5];
assign h2f_lw_WDATA[6] = hps2fpga_light_weight_WDATA_bus[6];
assign h2f_lw_WDATA[7] = hps2fpga_light_weight_WDATA_bus[7];
assign h2f_lw_WDATA[8] = hps2fpga_light_weight_WDATA_bus[8];
assign h2f_lw_WDATA[9] = hps2fpga_light_weight_WDATA_bus[9];
assign h2f_lw_WDATA[10] = hps2fpga_light_weight_WDATA_bus[10];
assign h2f_lw_WDATA[11] = hps2fpga_light_weight_WDATA_bus[11];
assign h2f_lw_WDATA[12] = hps2fpga_light_weight_WDATA_bus[12];
assign h2f_lw_WDATA[13] = hps2fpga_light_weight_WDATA_bus[13];
assign h2f_lw_WDATA[14] = hps2fpga_light_weight_WDATA_bus[14];
assign h2f_lw_WDATA[15] = hps2fpga_light_weight_WDATA_bus[15];
assign h2f_lw_WDATA[16] = hps2fpga_light_weight_WDATA_bus[16];
assign h2f_lw_WDATA[17] = hps2fpga_light_weight_WDATA_bus[17];
assign h2f_lw_WDATA[18] = hps2fpga_light_weight_WDATA_bus[18];
assign h2f_lw_WDATA[19] = hps2fpga_light_weight_WDATA_bus[19];
assign h2f_lw_WDATA[20] = hps2fpga_light_weight_WDATA_bus[20];
assign h2f_lw_WDATA[21] = hps2fpga_light_weight_WDATA_bus[21];
assign h2f_lw_WDATA[22] = hps2fpga_light_weight_WDATA_bus[22];
assign h2f_lw_WDATA[23] = hps2fpga_light_weight_WDATA_bus[23];
assign h2f_lw_WDATA[24] = hps2fpga_light_weight_WDATA_bus[24];
assign h2f_lw_WDATA[25] = hps2fpga_light_weight_WDATA_bus[25];
assign h2f_lw_WDATA[26] = hps2fpga_light_weight_WDATA_bus[26];
assign h2f_lw_WDATA[27] = hps2fpga_light_weight_WDATA_bus[27];
assign h2f_lw_WDATA[28] = hps2fpga_light_weight_WDATA_bus[28];
assign h2f_lw_WDATA[29] = hps2fpga_light_weight_WDATA_bus[29];
assign h2f_lw_WDATA[30] = hps2fpga_light_weight_WDATA_bus[30];
assign h2f_lw_WDATA[31] = hps2fpga_light_weight_WDATA_bus[31];

assign h2f_lw_WSTRB[0] = hps2fpga_light_weight_WSTRB_bus[0];
assign h2f_lw_WSTRB[1] = hps2fpga_light_weight_WSTRB_bus[1];
assign h2f_lw_WSTRB[2] = hps2fpga_light_weight_WSTRB_bus[2];
assign h2f_lw_WSTRB[3] = hps2fpga_light_weight_WSTRB_bus[3];

cyclonev_hps_interface_clocks_resets clocks_resets(
	.f2h_cold_rst_req_n(vcc),
	.f2h_dbg_rst_req_n(vcc),
	.f2h_pending_rst_ack(vcc),
	.f2h_periph_ref_clk(gnd),
	.f2h_sdram_ref_clk(gnd),
	.f2h_warm_rst_req_n(vcc),
	.ptp_ref_clk(gnd),
	.h2f_cold_rst_n(\clocks_resets~h2f_cold_rst_n ),
	.h2f_pending_rst_req_n(),
	.h2f_rst_n(h2f_rst_n[0]),
	.h2f_user0_clk(),
	.h2f_user1_clk(),
	.h2f_user2_clk());
defparam clocks_resets.h2f_user0_clk_freq = 100;
defparam clocks_resets.h2f_user1_clk_freq = 100;
defparam clocks_resets.h2f_user2_clk_freq = 100;

cyclonev_hps_interface_hps2fpga_light_weight hps2fpga_light_weight(
	.arready(h2f_lw_ARREADY[0]),
	.awready(h2f_lw_AWREADY[0]),
	.bvalid(h2f_lw_BVALID[0]),
	.clk(f2h_axi_clk[0]),
	.rlast(h2f_lw_RLAST[0]),
	.rvalid(h2f_lw_RVALID[0]),
	.wready(h2f_lw_WREADY[0]),
	.bid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.bresp({gnd,gnd}),
	.rdata({h2f_lw_RDATA[31],h2f_lw_RDATA[30],h2f_lw_RDATA[29],h2f_lw_RDATA[28],h2f_lw_RDATA[27],h2f_lw_RDATA[26],h2f_lw_RDATA[25],h2f_lw_RDATA[24],h2f_lw_RDATA[23],h2f_lw_RDATA[22],h2f_lw_RDATA[21],h2f_lw_RDATA[20],h2f_lw_RDATA[19],h2f_lw_RDATA[18],h2f_lw_RDATA[17],h2f_lw_RDATA[16],h2f_lw_RDATA[15],h2f_lw_RDATA[14],h2f_lw_RDATA[13],h2f_lw_RDATA[12],h2f_lw_RDATA[11],
h2f_lw_RDATA[10],h2f_lw_RDATA[9],h2f_lw_RDATA[8],h2f_lw_RDATA[7],h2f_lw_RDATA[6],h2f_lw_RDATA[5],h2f_lw_RDATA[4],h2f_lw_RDATA[3],h2f_lw_RDATA[2],h2f_lw_RDATA[1],h2f_lw_RDATA[0]}),
	.rid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_lw_ARVALID[0]),
	.awvalid(h2f_lw_AWVALID[0]),
	.bready(h2f_lw_BREADY[0]),
	.rready(h2f_lw_RREADY[0]),
	.wlast(h2f_lw_WLAST[0]),
	.wvalid(h2f_lw_WVALID[0]),
	.araddr(hps2fpga_light_weight_ARADDR_bus),
	.arburst(hps2fpga_light_weight_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_light_weight_ARID_bus),
	.arlen(hps2fpga_light_weight_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_light_weight_ARSIZE_bus),
	.awaddr(hps2fpga_light_weight_AWADDR_bus),
	.awburst(hps2fpga_light_weight_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_light_weight_AWID_bus),
	.awlen(hps2fpga_light_weight_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_light_weight_AWSIZE_bus),
	.wdata(hps2fpga_light_weight_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_light_weight_WSTRB_bus));

cyclonev_hps_interface_dbg_apb debug_apb(
	.p_slv_err(gnd),
	.p_ready(gnd),
	.p_clk(gnd),
	.p_clk_en(gnd),
	.dbg_apb_disable(gnd),
	.p_rdata(32'b00000000000000000000000000000000),
	.p_addr_31(\debug_apb~O_P_ADDR_31 ),
	.p_write(),
	.p_sel(),
	.p_enable(),
	.p_reset_n(),
	.p_addr(),
	.p_wdata());
defparam debug_apb.dummy_param = 256;

cyclonev_hps_interface_tpiu_trace tpiu(
	.traceclk_ctl(vcc),
	.traceclkin(gnd),
	.traceclk(),
	.trace_data(tpiu_TRACE_DATA_bus));

cyclonev_hps_interface_boot_from_fpga boot_from_fpga(
	.boot_from_fpga_on_failure(gnd),
	.boot_from_fpga_ready(gnd),
	.bsel_en(gnd),
	.csel_en(gnd),
	.bsel({gnd,gnd,vcc}),
	.csel({gnd,vcc}),
	.fake_dout(\boot_from_fpga~fake_dout ));

cyclonev_hps_interface_fpga2hps fpga2hps(
	.arvalid(gnd),
	.awvalid(gnd),
	.bready(gnd),
	.clk(f2h_axi_clk[0]),
	.rready(gnd),
	.wlast(gnd),
	.wvalid(gnd),
	.araddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arburst({gnd,gnd}),
	.arcache({gnd,gnd,gnd,gnd}),
	.arid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arlen({gnd,gnd,gnd,gnd}),
	.arlock({gnd,gnd}),
	.arprot({gnd,gnd,gnd}),
	.arsize({gnd,gnd,gnd}),
	.aruser({gnd,gnd,gnd,gnd,gnd}),
	.awaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awburst({gnd,gnd}),
	.awcache({gnd,gnd,gnd,gnd}),
	.awid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awlen({gnd,gnd,gnd,gnd}),
	.awlock({gnd,gnd}),
	.awprot({gnd,gnd,gnd}),
	.awsize({gnd,gnd,gnd}),
	.awuser({gnd,gnd,gnd,gnd,gnd}),
	.port_size_config({gnd,vcc}),
	.wdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wstrb({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arready(\f2h_ARREADY[0] ),
	.awready(),
	.bvalid(),
	.rlast(),
	.rvalid(),
	.wready(),
	.bid(),
	.bresp(),
	.rdata(),
	.rid(),
	.rresp());
defparam fpga2hps.data_width = 32;

cyclonev_hps_interface_hps2fpga hps2fpga(
	.arready(gnd),
	.awready(gnd),
	.bvalid(gnd),
	.clk(f2h_axi_clk[0]),
	.rlast(gnd),
	.rvalid(gnd),
	.wready(gnd),
	.bid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.bresp({gnd,gnd}),
	.port_size_config({vcc,gnd}),
	.rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rresp({gnd,gnd}),
	.arvalid(),
	.awvalid(),
	.bready(),
	.rready(),
	.wlast(),
	.wvalid(),
	.araddr(hps2fpga_ARADDR_bus),
	.arburst(),
	.arcache(),
	.arid(),
	.arlen(),
	.arlock(),
	.arprot(),
	.arsize(),
	.awaddr(),
	.awburst(),
	.awcache(),
	.awid(),
	.awlen(),
	.awlock(),
	.awprot(),
	.awsize(),
	.wdata(),
	.wid(),
	.wstrb());
defparam hps2fpga.data_width = 32;

cyclonev_hps_interface_fpga2sdram f2sdram(
	.cmd_port_clk_0(gnd),
	.cmd_port_clk_1(gnd),
	.cmd_port_clk_2(gnd),
	.cmd_port_clk_3(gnd),
	.cmd_port_clk_4(gnd),
	.cmd_port_clk_5(gnd),
	.cmd_valid_0(gnd),
	.cmd_valid_1(gnd),
	.cmd_valid_2(gnd),
	.cmd_valid_3(gnd),
	.cmd_valid_4(gnd),
	.cmd_valid_5(gnd),
	.rd_clk_0(gnd),
	.rd_clk_1(gnd),
	.rd_clk_2(gnd),
	.rd_clk_3(gnd),
	.rd_ready_0(gnd),
	.rd_ready_1(gnd),
	.rd_ready_2(gnd),
	.rd_ready_3(gnd),
	.wr_clk_0(gnd),
	.wr_clk_1(gnd),
	.wr_clk_2(gnd),
	.wr_clk_3(gnd),
	.wr_valid_0(gnd),
	.wr_valid_1(gnd),
	.wr_valid_2(gnd),
	.wr_valid_3(gnd),
	.wrack_ready_0(gnd),
	.wrack_ready_1(gnd),
	.wrack_ready_2(gnd),
	.wrack_ready_3(gnd),
	.wrack_ready_4(gnd),
	.wrack_ready_5(gnd),
	.cfg_axi_mm_select({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_rfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_type({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_wfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_port_width({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_rfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_wfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_data_0(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_1(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_2(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_3(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_4(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_5(60'b000000000000000000000000000000000000000000000000000000000000),
	.wr_data_0(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_1(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_2(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_3(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.cmd_ready_0(),
	.cmd_ready_1(),
	.cmd_ready_2(),
	.cmd_ready_3(),
	.cmd_ready_4(),
	.cmd_ready_5(),
	.rd_valid_0(),
	.rd_valid_1(),
	.rd_valid_2(),
	.rd_valid_3(),
	.wr_ready_0(),
	.wr_ready_1(),
	.wr_ready_2(),
	.wr_ready_3(),
	.wrack_valid_0(),
	.wrack_valid_1(),
	.wrack_valid_2(),
	.wrack_valid_3(),
	.wrack_valid_4(),
	.wrack_valid_5(),
	.bonding_out_1(f2sdram_BONDING_OUT_1_bus),
	.bonding_out_2(),
	.rd_data_0(),
	.rd_data_1(),
	.rd_data_2(),
	.rd_data_3(),
	.wrack_data_0(),
	.wrack_data_1(),
	.wrack_data_2(),
	.wrack_data_3(),
	.wrack_data_4(),
	.wrack_data_5());

cyclonev_hps_interface_interrupts interrupts(
	.irq({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.fake_dout(\interrupts~fake_dout ),
	.h2f_can0_irq(),
	.h2f_can1_irq(),
	.h2f_clkmgr_irq(),
	.h2f_cti_irq0_n(),
	.h2f_cti_irq1_n(),
	.h2f_dma_abort_irq(),
	.h2f_dma_irq0(),
	.h2f_dma_irq1(),
	.h2f_dma_irq2(),
	.h2f_dma_irq3(),
	.h2f_dma_irq4(),
	.h2f_dma_irq5(),
	.h2f_dma_irq6(),
	.h2f_dma_irq7(),
	.h2f_emac0_irq(),
	.h2f_emac1_irq(),
	.h2f_fpga_man_irq(),
	.h2f_gpio0_irq(),
	.h2f_gpio1_irq(),
	.h2f_gpio2_irq(),
	.h2f_i2c0_irq(),
	.h2f_i2c1_irq(),
	.h2f_i2c_emac0_irq(),
	.h2f_i2c_emac1_irq(),
	.h2f_l4sp0_irq(),
	.h2f_l4sp1_irq(),
	.h2f_mpuwakeup_irq(),
	.h2f_nand_irq(),
	.h2f_osc0_irq(),
	.h2f_osc1_irq(),
	.h2f_qspi_irq(),
	.h2f_sdmmc_irq(),
	.h2f_spi0_irq(),
	.h2f_spi1_irq(),
	.h2f_spi2_irq(),
	.h2f_spi3_irq(),
	.h2f_uart0_irq(),
	.h2f_uart1_irq(),
	.h2f_usb0_irq(),
	.h2f_usb1_irq(),
	.h2f_wdog0_irq(),
	.h2f_wdog1_irq());

endmodule

module system_system_hps_0_hps_io (
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim1_inst,
	spim1_inst1,
	intermediate_36,
	intermediate_37,
	uart0_inst,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	uart0_inst;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_system_hps_0_hps_io_border border(
	.hps_io_emac1_inst_TX_CLK({emac1_inst}),
	.hps_io_emac1_inst_TX_CTL({emac1_inst1}),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.hps_io_emac1_inst_MDC({emac1_inst2}),
	.hps_io_emac1_inst_TXD0({emac1_inst3}),
	.hps_io_emac1_inst_TXD1({emac1_inst4}),
	.hps_io_emac1_inst_TXD2({emac1_inst5}),
	.hps_io_emac1_inst_TXD3({emac1_inst6}),
	.hps_io_qspi_inst_CLK({qspi_inst}),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.hps_io_qspi_inst_SS0({qspi_inst1}),
	.hps_io_sdio_inst_CLK({sdio_inst}),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.hps_io_usb1_inst_STP({usb1_inst}),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.hps_io_spim1_inst_CLK({spim1_inst}),
	.hps_io_spim1_inst_SS0({spim1_inst1}),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.hps_io_uart0_inst_TX({uart0_inst}),
	.intermediate_39(intermediate_39),
	.intermediate_38(intermediate_38),
	.intermediate_41(intermediate_41),
	.intermediate_40(intermediate_40),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_i2c0_inst_SDA_0(hps_io_i2c0_inst_SDA_0),
	.hps_io_i2c0_inst_SCL_0(hps_io_i2c0_inst_SCL_0),
	.hps_io_i2c1_inst_SDA_0(hps_io_i2c1_inst_SDA_0),
	.hps_io_i2c1_inst_SCL_0(hps_io_i2c1_inst_SCL_0),
	.hps_io_emac1_inst_RXD0({hps_io_hps_io_emac1_inst_RXD0}),
	.hps_io_emac1_inst_RXD1({hps_io_hps_io_emac1_inst_RXD1}),
	.hps_io_emac1_inst_RXD2({hps_io_hps_io_emac1_inst_RXD2}),
	.hps_io_emac1_inst_RXD3({hps_io_hps_io_emac1_inst_RXD3}),
	.hps_io_emac1_inst_RX_CLK({hps_io_hps_io_emac1_inst_RX_CLK}),
	.hps_io_emac1_inst_RX_CTL({hps_io_hps_io_emac1_inst_RX_CTL}),
	.hps_io_spim1_inst_MISO({hps_io_hps_io_spim1_inst_MISO}),
	.hps_io_uart0_inst_RX({hps_io_hps_io_uart0_inst_RX}),
	.hps_io_usb1_inst_CLK({hps_io_hps_io_usb1_inst_CLK}),
	.hps_io_usb1_inst_DIR({hps_io_hps_io_usb1_inst_DIR}),
	.hps_io_usb1_inst_NXT({hps_io_hps_io_usb1_inst_NXT}),
	.memory_oct_rzqin(memory_oct_rzqin));

endmodule

module system_system_hps_0_hps_io_border (
	hps_io_emac1_inst_TX_CLK,
	hps_io_emac1_inst_TX_CTL,
	intermediate_0,
	intermediate_1,
	hps_io_emac1_inst_MDC,
	hps_io_emac1_inst_TXD0,
	hps_io_emac1_inst_TXD1,
	hps_io_emac1_inst_TXD2,
	hps_io_emac1_inst_TXD3,
	hps_io_qspi_inst_CLK,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	hps_io_qspi_inst_SS0,
	hps_io_sdio_inst_CLK,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	hps_io_usb1_inst_STP,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	hps_io_spim1_inst_CLK,
	hps_io_spim1_inst_SS0,
	intermediate_36,
	intermediate_37,
	hps_io_uart0_inst_TX,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_emac1_inst_RXD0,
	hps_io_emac1_inst_RXD1,
	hps_io_emac1_inst_RXD2,
	hps_io_emac1_inst_RXD3,
	hps_io_emac1_inst_RX_CLK,
	hps_io_emac1_inst_RX_CTL,
	hps_io_spim1_inst_MISO,
	hps_io_uart0_inst_RX,
	hps_io_usb1_inst_CLK,
	hps_io_usb1_inst_DIR,
	hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[0:0] hps_io_emac1_inst_TX_CLK;
output 	[0:0] hps_io_emac1_inst_TX_CTL;
output 	intermediate_0;
output 	intermediate_1;
output 	[0:0] hps_io_emac1_inst_MDC;
output 	[0:0] hps_io_emac1_inst_TXD0;
output 	[0:0] hps_io_emac1_inst_TXD1;
output 	[0:0] hps_io_emac1_inst_TXD2;
output 	[0:0] hps_io_emac1_inst_TXD3;
output 	[0:0] hps_io_qspi_inst_CLK;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	[0:0] hps_io_qspi_inst_SS0;
output 	[0:0] hps_io_sdio_inst_CLK;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	[0:0] hps_io_usb1_inst_STP;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	[0:0] hps_io_spim1_inst_CLK;
output 	[0:0] hps_io_spim1_inst_SS0;
output 	intermediate_36;
output 	intermediate_37;
output 	[0:0] hps_io_uart0_inst_TX;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	[0:0] hps_io_emac1_inst_RXD0;
input 	[0:0] hps_io_emac1_inst_RXD1;
input 	[0:0] hps_io_emac1_inst_RXD2;
input 	[0:0] hps_io_emac1_inst_RXD3;
input 	[0:0] hps_io_emac1_inst_RX_CLK;
input 	[0:0] hps_io_emac1_inst_RX_CTL;
input 	[0:0] hps_io_spim1_inst_MISO;
input 	[0:0] hps_io_uart0_inst_RX;
input 	[0:0] hps_io_usb1_inst_CLK;
input 	[0:0] hps_io_usb1_inst_DIR;
input 	[0:0] hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdio_inst~O_SDMMC_PWR_EN ;
wire \uart0_inst~UARTRTSN ;
wire \~GND~combout ;

wire [3:0] emac1_inst_EMAC_PHY_TXD_bus;
wire [3:0] qspi_inst_QSPI_SS_N_bus;
wire [3:0] qspi_inst_QSPI_MO_EN_N_bus;
wire [7:0] sdio_inst_SDMMC_DATA_OE_bus;
wire [7:0] sdio_inst_SDMMC_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_OE_bus;

assign hps_io_emac1_inst_TXD0[0] = emac1_inst_EMAC_PHY_TXD_bus[0];
assign hps_io_emac1_inst_TXD1[0] = emac1_inst_EMAC_PHY_TXD_bus[1];
assign hps_io_emac1_inst_TXD2[0] = emac1_inst_EMAC_PHY_TXD_bus[2];
assign hps_io_emac1_inst_TXD3[0] = emac1_inst_EMAC_PHY_TXD_bus[3];

assign hps_io_qspi_inst_SS0[0] = qspi_inst_QSPI_SS_N_bus[0];

assign intermediate_3 = qspi_inst_QSPI_MO_EN_N_bus[0];
assign intermediate_5 = qspi_inst_QSPI_MO_EN_N_bus[1];
assign intermediate_7 = qspi_inst_QSPI_MO_EN_N_bus[2];
assign intermediate_9 = qspi_inst_QSPI_MO_EN_N_bus[3];

assign intermediate_13 = sdio_inst_SDMMC_DATA_OE_bus[0];
assign intermediate_15 = sdio_inst_SDMMC_DATA_OE_bus[1];
assign intermediate_17 = sdio_inst_SDMMC_DATA_OE_bus[2];
assign intermediate_19 = sdio_inst_SDMMC_DATA_OE_bus[3];

assign intermediate_12 = sdio_inst_SDMMC_DATA_O_bus[0];
assign intermediate_14 = sdio_inst_SDMMC_DATA_O_bus[1];
assign intermediate_16 = sdio_inst_SDMMC_DATA_O_bus[2];
assign intermediate_18 = sdio_inst_SDMMC_DATA_O_bus[3];

assign intermediate_20 = usb1_inst_USB_ULPI_DATA_O_bus[0];
assign intermediate_22 = usb1_inst_USB_ULPI_DATA_O_bus[1];
assign intermediate_24 = usb1_inst_USB_ULPI_DATA_O_bus[2];
assign intermediate_26 = usb1_inst_USB_ULPI_DATA_O_bus[3];
assign intermediate_28 = usb1_inst_USB_ULPI_DATA_O_bus[4];
assign intermediate_30 = usb1_inst_USB_ULPI_DATA_O_bus[5];
assign intermediate_32 = usb1_inst_USB_ULPI_DATA_O_bus[6];
assign intermediate_34 = usb1_inst_USB_ULPI_DATA_O_bus[7];

assign intermediate_21 = usb1_inst_USB_ULPI_DATA_OE_bus[0];
assign intermediate_23 = usb1_inst_USB_ULPI_DATA_OE_bus[1];
assign intermediate_25 = usb1_inst_USB_ULPI_DATA_OE_bus[2];
assign intermediate_27 = usb1_inst_USB_ULPI_DATA_OE_bus[3];
assign intermediate_29 = usb1_inst_USB_ULPI_DATA_OE_bus[4];
assign intermediate_31 = usb1_inst_USB_ULPI_DATA_OE_bus[5];
assign intermediate_33 = usb1_inst_USB_ULPI_DATA_OE_bus[6];
assign intermediate_35 = usb1_inst_USB_ULPI_DATA_OE_bus[7];

system_hps_sdram hps_sdram_inst(
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.GND_port(\~GND~combout ),
	.memory_oct_rzqin(memory_oct_rzqin));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_hps_peripheral_emac emac1_inst(
	.emac_clk_rx(hps_io_emac1_inst_RX_CLK[0]),
	.emac_phy_rxdv(hps_io_emac1_inst_RX_CTL[0]),
	.emac_gmii_mdo_i(hps_io_emac1_inst_MDIO_0),
	.emac_phy_rxd({hps_io_emac1_inst_RXD3[0],hps_io_emac1_inst_RXD2[0],hps_io_emac1_inst_RXD1[0],hps_io_emac1_inst_RXD0[0]}),
	.emac_clk_tx(hps_io_emac1_inst_TX_CLK[0]),
	.emac_phy_tx_oe(hps_io_emac1_inst_TX_CTL[0]),
	.emac_gmii_mdo_o(intermediate_0),
	.emac_gmii_mdo_oe(intermediate_1),
	.emac_gmii_mdc(hps_io_emac1_inst_MDC[0]),
	.emac_phy_txd(emac1_inst_EMAC_PHY_TXD_bus));
defparam emac1_inst.dummy_param = 256;

cyclonev_hps_peripheral_qspi qspi_inst(
	.qspi_mi0(hps_io_qspi_inst_IO0_0),
	.qspi_mi1(hps_io_qspi_inst_IO1_0),
	.qspi_mi2(hps_io_qspi_inst_IO2_0),
	.qspi_mi3(hps_io_qspi_inst_IO3_0),
	.qspi_sclk(hps_io_qspi_inst_CLK[0]),
	.qspi_mo0(intermediate_2),
	.qspi_mo1(intermediate_4),
	.qspi_mo2(intermediate_6),
	.qspi_mo3(intermediate_8),
	.qspi_mo_en_n(qspi_inst_QSPI_MO_EN_N_bus),
	.qspi_ss_n(qspi_inst_QSPI_SS_N_bus));
defparam qspi_inst.dummy_param = 256;

cyclonev_hps_peripheral_sdmmc sdio_inst(
	.sdmmc_fb_clk(gnd),
	.sdmmc_cmd_i(hps_io_sdio_inst_CMD_0),
	.sdmmc_data_i({gnd,gnd,gnd,gnd,hps_io_sdio_inst_D3_0,hps_io_sdio_inst_D2_0,hps_io_sdio_inst_D1_0,hps_io_sdio_inst_D0_0}),
	.sdmmc_pwr_en(\sdio_inst~O_SDMMC_PWR_EN ),
	.sdmmc_cclk(hps_io_sdio_inst_CLK[0]),
	.sdmmc_cmd_o(intermediate_10),
	.sdmmc_cmd_oe(intermediate_11),
	.sdmmc_data_o(sdio_inst_SDMMC_DATA_O_bus),
	.sdmmc_data_oe(sdio_inst_SDMMC_DATA_OE_bus));
defparam sdio_inst.dummy_param = 256;

cyclonev_hps_peripheral_usb usb1_inst(
	.usb_ulpi_clk(hps_io_usb1_inst_CLK[0]),
	.usb_ulpi_dir(hps_io_usb1_inst_DIR[0]),
	.usb_ulpi_nxt(hps_io_usb1_inst_NXT[0]),
	.usb_ulpi_data_i({hps_io_usb1_inst_D7_0,hps_io_usb1_inst_D6_0,hps_io_usb1_inst_D5_0,hps_io_usb1_inst_D4_0,hps_io_usb1_inst_D3_0,hps_io_usb1_inst_D2_0,hps_io_usb1_inst_D1_0,hps_io_usb1_inst_D0_0}),
	.usb_ulpi_stp(hps_io_usb1_inst_STP[0]),
	.usb_ulpi_data_o(usb1_inst_USB_ULPI_DATA_O_bus),
	.usb_ulpi_data_oe(usb1_inst_USB_ULPI_DATA_OE_bus));
defparam usb1_inst.dummy_param = 256;

cyclonev_hps_peripheral_spi_master spim1_inst(
	.spi_master_rxd(hps_io_spim1_inst_MISO[0]),
	.spi_master_sclk(hps_io_spim1_inst_CLK[0]),
	.spi_master_ss_0_n(hps_io_spim1_inst_SS0[0]),
	.spi_master_ss_1_n(),
	.spi_master_txd(intermediate_36),
	.spi_master_ssi_oe_n(intermediate_37));
defparam spim1_inst.dummy_param = 256;

cyclonev_hps_peripheral_uart uart0_inst(
	.uart_cts_n(gnd),
	.uart_rxd(hps_io_uart0_inst_RX[0]),
	.uart_rts_n(\uart0_inst~UARTRTSN ),
	.uart_txd(hps_io_uart0_inst_TX[0]));
defparam uart0_inst.dummy_param = 256;

cyclonev_hps_peripheral_i2c i2c0_inst(
	.i2c_clk(hps_io_i2c0_inst_SCL_0),
	.i2c_data(hps_io_i2c0_inst_SDA_0),
	.i2c_clk_oe(intermediate_39),
	.i2c_data_oe(intermediate_38));
defparam i2c0_inst.dummy_param = 256;

cyclonev_hps_peripheral_i2c i2c1_inst(
	.i2c_clk(hps_io_i2c1_inst_SCL_0),
	.i2c_data(hps_io_i2c1_inst_SDA_0),
	.i2c_clk_oe(intermediate_41),
	.i2c_data_oe(intermediate_40));
defparam i2c1_inst.dummy_param = 256;

endmodule

module system_hps_sdram (
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	GND_port,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	GND_port;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pll|afi_clk ;
wire \pll|pll_write_clk ;
wire \p0|umemphy|afi_cal_fail ;
wire \p0|umemphy|afi_cal_success ;
wire \p0|umemphy|afi_rdata_valid[0] ;
wire \p0|umemphy|ctl_reset_n ;
wire \p0|umemphy|afi_rdata[0] ;
wire \p0|umemphy|afi_rdata[1] ;
wire \p0|umemphy|afi_rdata[2] ;
wire \p0|umemphy|afi_rdata[3] ;
wire \p0|umemphy|afi_rdata[4] ;
wire \p0|umemphy|afi_rdata[5] ;
wire \p0|umemphy|afi_rdata[6] ;
wire \p0|umemphy|afi_rdata[7] ;
wire \p0|umemphy|afi_rdata[8] ;
wire \p0|umemphy|afi_rdata[9] ;
wire \p0|umemphy|afi_rdata[10] ;
wire \p0|umemphy|afi_rdata[11] ;
wire \p0|umemphy|afi_rdata[12] ;
wire \p0|umemphy|afi_rdata[13] ;
wire \p0|umemphy|afi_rdata[14] ;
wire \p0|umemphy|afi_rdata[15] ;
wire \p0|umemphy|afi_rdata[16] ;
wire \p0|umemphy|afi_rdata[17] ;
wire \p0|umemphy|afi_rdata[18] ;
wire \p0|umemphy|afi_rdata[19] ;
wire \p0|umemphy|afi_rdata[20] ;
wire \p0|umemphy|afi_rdata[21] ;
wire \p0|umemphy|afi_rdata[22] ;
wire \p0|umemphy|afi_rdata[23] ;
wire \p0|umemphy|afi_rdata[24] ;
wire \p0|umemphy|afi_rdata[25] ;
wire \p0|umemphy|afi_rdata[26] ;
wire \p0|umemphy|afi_rdata[27] ;
wire \p0|umemphy|afi_rdata[28] ;
wire \p0|umemphy|afi_rdata[29] ;
wire \p0|umemphy|afi_rdata[30] ;
wire \p0|umemphy|afi_rdata[31] ;
wire \p0|umemphy|afi_rdata[32] ;
wire \p0|umemphy|afi_rdata[33] ;
wire \p0|umemphy|afi_rdata[34] ;
wire \p0|umemphy|afi_rdata[35] ;
wire \p0|umemphy|afi_rdata[36] ;
wire \p0|umemphy|afi_rdata[37] ;
wire \p0|umemphy|afi_rdata[38] ;
wire \p0|umemphy|afi_rdata[39] ;
wire \p0|umemphy|afi_rdata[40] ;
wire \p0|umemphy|afi_rdata[41] ;
wire \p0|umemphy|afi_rdata[42] ;
wire \p0|umemphy|afi_rdata[43] ;
wire \p0|umemphy|afi_rdata[44] ;
wire \p0|umemphy|afi_rdata[45] ;
wire \p0|umemphy|afi_rdata[46] ;
wire \p0|umemphy|afi_rdata[47] ;
wire \p0|umemphy|afi_rdata[48] ;
wire \p0|umemphy|afi_rdata[49] ;
wire \p0|umemphy|afi_rdata[50] ;
wire \p0|umemphy|afi_rdata[51] ;
wire \p0|umemphy|afi_rdata[52] ;
wire \p0|umemphy|afi_rdata[53] ;
wire \p0|umemphy|afi_rdata[54] ;
wire \p0|umemphy|afi_rdata[55] ;
wire \p0|umemphy|afi_rdata[56] ;
wire \p0|umemphy|afi_rdata[57] ;
wire \p0|umemphy|afi_rdata[58] ;
wire \p0|umemphy|afi_rdata[59] ;
wire \p0|umemphy|afi_rdata[60] ;
wire \p0|umemphy|afi_rdata[61] ;
wire \p0|umemphy|afi_rdata[62] ;
wire \p0|umemphy|afi_rdata[63] ;
wire \p0|umemphy|afi_rdata[64] ;
wire \p0|umemphy|afi_rdata[65] ;
wire \p0|umemphy|afi_rdata[66] ;
wire \p0|umemphy|afi_rdata[67] ;
wire \p0|umemphy|afi_rdata[68] ;
wire \p0|umemphy|afi_rdata[69] ;
wire \p0|umemphy|afi_rdata[70] ;
wire \p0|umemphy|afi_rdata[71] ;
wire \p0|umemphy|afi_rdata[72] ;
wire \p0|umemphy|afi_rdata[73] ;
wire \p0|umemphy|afi_rdata[74] ;
wire \p0|umemphy|afi_rdata[75] ;
wire \p0|umemphy|afi_rdata[76] ;
wire \p0|umemphy|afi_rdata[77] ;
wire \p0|umemphy|afi_rdata[78] ;
wire \p0|umemphy|afi_rdata[79] ;
wire \p0|umemphy|afi_wlat[0] ;
wire \p0|umemphy|afi_wlat[1] ;
wire \p0|umemphy|afi_wlat[2] ;
wire \p0|umemphy|afi_wlat[3] ;
wire \c0|afi_cas_n[0] ;
wire \c0|afi_ras_n[0] ;
wire \c0|afi_rst_n[0] ;
wire \c0|afi_we_n[0] ;
wire \c0|afi_addr[0] ;
wire \c0|afi_addr[1] ;
wire \c0|afi_addr[2] ;
wire \c0|afi_addr[3] ;
wire \c0|afi_addr[4] ;
wire \c0|afi_addr[5] ;
wire \c0|afi_addr[6] ;
wire \c0|afi_addr[7] ;
wire \c0|afi_addr[8] ;
wire \c0|afi_addr[9] ;
wire \c0|afi_addr[10] ;
wire \c0|afi_addr[11] ;
wire \c0|afi_addr[12] ;
wire \c0|afi_addr[13] ;
wire \c0|afi_addr[14] ;
wire \c0|afi_addr[15] ;
wire \c0|afi_addr[16] ;
wire \c0|afi_addr[17] ;
wire \c0|afi_addr[18] ;
wire \c0|afi_addr[19] ;
wire \c0|afi_ba[0] ;
wire \c0|afi_ba[1] ;
wire \c0|afi_ba[2] ;
wire \c0|afi_cke[0] ;
wire \c0|afi_cke[1] ;
wire \c0|afi_cs_n[0] ;
wire \c0|afi_cs_n[1] ;
wire \c0|afi_dm_int[0] ;
wire \c0|afi_dm_int[1] ;
wire \c0|afi_dm_int[2] ;
wire \c0|afi_dm_int[3] ;
wire \c0|afi_dm_int[4] ;
wire \c0|afi_dm_int[5] ;
wire \c0|afi_dm_int[6] ;
wire \c0|afi_dm_int[7] ;
wire \c0|afi_dm_int[8] ;
wire \c0|afi_dm_int[9] ;
wire \c0|afi_dqs_burst[0] ;
wire \c0|afi_dqs_burst[1] ;
wire \c0|afi_dqs_burst[2] ;
wire \c0|afi_dqs_burst[3] ;
wire \c0|afi_dqs_burst[4] ;
wire \c0|afi_odt[0] ;
wire \c0|afi_odt[1] ;
wire \c0|afi_rdata_en[0] ;
wire \c0|afi_rdata_en[1] ;
wire \c0|afi_rdata_en[2] ;
wire \c0|afi_rdata_en[3] ;
wire \c0|afi_rdata_en[4] ;
wire \c0|afi_rdata_en_full[0] ;
wire \c0|afi_rdata_en_full[1] ;
wire \c0|afi_rdata_en_full[2] ;
wire \c0|afi_rdata_en_full[3] ;
wire \c0|afi_rdata_en_full[4] ;
wire \c0|afi_wdata_int[0] ;
wire \c0|afi_wdata_int[1] ;
wire \c0|afi_wdata_int[2] ;
wire \c0|afi_wdata_int[3] ;
wire \c0|afi_wdata_int[4] ;
wire \c0|afi_wdata_int[5] ;
wire \c0|afi_wdata_int[6] ;
wire \c0|afi_wdata_int[7] ;
wire \c0|afi_wdata_int[8] ;
wire \c0|afi_wdata_int[9] ;
wire \c0|afi_wdata_int[10] ;
wire \c0|afi_wdata_int[11] ;
wire \c0|afi_wdata_int[12] ;
wire \c0|afi_wdata_int[13] ;
wire \c0|afi_wdata_int[14] ;
wire \c0|afi_wdata_int[15] ;
wire \c0|afi_wdata_int[16] ;
wire \c0|afi_wdata_int[17] ;
wire \c0|afi_wdata_int[18] ;
wire \c0|afi_wdata_int[19] ;
wire \c0|afi_wdata_int[20] ;
wire \c0|afi_wdata_int[21] ;
wire \c0|afi_wdata_int[22] ;
wire \c0|afi_wdata_int[23] ;
wire \c0|afi_wdata_int[24] ;
wire \c0|afi_wdata_int[25] ;
wire \c0|afi_wdata_int[26] ;
wire \c0|afi_wdata_int[27] ;
wire \c0|afi_wdata_int[28] ;
wire \c0|afi_wdata_int[29] ;
wire \c0|afi_wdata_int[30] ;
wire \c0|afi_wdata_int[31] ;
wire \c0|afi_wdata_int[32] ;
wire \c0|afi_wdata_int[33] ;
wire \c0|afi_wdata_int[34] ;
wire \c0|afi_wdata_int[35] ;
wire \c0|afi_wdata_int[36] ;
wire \c0|afi_wdata_int[37] ;
wire \c0|afi_wdata_int[38] ;
wire \c0|afi_wdata_int[39] ;
wire \c0|afi_wdata_int[40] ;
wire \c0|afi_wdata_int[41] ;
wire \c0|afi_wdata_int[42] ;
wire \c0|afi_wdata_int[43] ;
wire \c0|afi_wdata_int[44] ;
wire \c0|afi_wdata_int[45] ;
wire \c0|afi_wdata_int[46] ;
wire \c0|afi_wdata_int[47] ;
wire \c0|afi_wdata_int[48] ;
wire \c0|afi_wdata_int[49] ;
wire \c0|afi_wdata_int[50] ;
wire \c0|afi_wdata_int[51] ;
wire \c0|afi_wdata_int[52] ;
wire \c0|afi_wdata_int[53] ;
wire \c0|afi_wdata_int[54] ;
wire \c0|afi_wdata_int[55] ;
wire \c0|afi_wdata_int[56] ;
wire \c0|afi_wdata_int[57] ;
wire \c0|afi_wdata_int[58] ;
wire \c0|afi_wdata_int[59] ;
wire \c0|afi_wdata_int[60] ;
wire \c0|afi_wdata_int[61] ;
wire \c0|afi_wdata_int[62] ;
wire \c0|afi_wdata_int[63] ;
wire \c0|afi_wdata_int[64] ;
wire \c0|afi_wdata_int[65] ;
wire \c0|afi_wdata_int[66] ;
wire \c0|afi_wdata_int[67] ;
wire \c0|afi_wdata_int[68] ;
wire \c0|afi_wdata_int[69] ;
wire \c0|afi_wdata_int[70] ;
wire \c0|afi_wdata_int[71] ;
wire \c0|afi_wdata_int[72] ;
wire \c0|afi_wdata_int[73] ;
wire \c0|afi_wdata_int[74] ;
wire \c0|afi_wdata_int[75] ;
wire \c0|afi_wdata_int[76] ;
wire \c0|afi_wdata_int[77] ;
wire \c0|afi_wdata_int[78] ;
wire \c0|afi_wdata_int[79] ;
wire \c0|afi_wdata_valid[0] ;
wire \c0|afi_wdata_valid[1] ;
wire \c0|afi_wdata_valid[2] ;
wire \c0|afi_wdata_valid[3] ;
wire \c0|afi_wdata_valid[4] ;
wire \c0|cfg_addlat_wire[0] ;
wire \c0|cfg_addlat_wire[1] ;
wire \c0|cfg_addlat_wire[2] ;
wire \c0|cfg_addlat_wire[3] ;
wire \c0|cfg_addlat_wire[4] ;
wire \c0|cfg_bankaddrwidth_wire[0] ;
wire \c0|cfg_bankaddrwidth_wire[1] ;
wire \c0|cfg_bankaddrwidth_wire[2] ;
wire \c0|cfg_caswrlat_wire[0] ;
wire \c0|cfg_caswrlat_wire[1] ;
wire \c0|cfg_caswrlat_wire[2] ;
wire \c0|cfg_caswrlat_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[0] ;
wire \c0|cfg_coladdrwidth_wire[1] ;
wire \c0|cfg_coladdrwidth_wire[2] ;
wire \c0|cfg_coladdrwidth_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[4] ;
wire \c0|cfg_csaddrwidth_wire[0] ;
wire \c0|cfg_csaddrwidth_wire[1] ;
wire \c0|cfg_csaddrwidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[0] ;
wire \c0|cfg_devicewidth_wire[1] ;
wire \c0|cfg_devicewidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[0] ;
wire \c0|cfg_interfacewidth_wire[1] ;
wire \c0|cfg_interfacewidth_wire[2] ;
wire \c0|cfg_interfacewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[4] ;
wire \c0|cfg_interfacewidth_wire[5] ;
wire \c0|cfg_interfacewidth_wire[6] ;
wire \c0|cfg_interfacewidth_wire[7] ;
wire \c0|cfg_rowaddrwidth_wire[0] ;
wire \c0|cfg_rowaddrwidth_wire[1] ;
wire \c0|cfg_rowaddrwidth_wire[2] ;
wire \c0|cfg_rowaddrwidth_wire[3] ;
wire \c0|cfg_rowaddrwidth_wire[4] ;
wire \c0|cfg_tcl_wire[0] ;
wire \c0|cfg_tcl_wire[1] ;
wire \c0|cfg_tcl_wire[2] ;
wire \c0|cfg_tcl_wire[3] ;
wire \c0|cfg_tcl_wire[4] ;
wire \c0|cfg_tmrd_wire[0] ;
wire \c0|cfg_tmrd_wire[1] ;
wire \c0|cfg_tmrd_wire[2] ;
wire \c0|cfg_tmrd_wire[3] ;
wire \c0|cfg_trefi_wire[0] ;
wire \c0|cfg_trefi_wire[1] ;
wire \c0|cfg_trefi_wire[2] ;
wire \c0|cfg_trefi_wire[3] ;
wire \c0|cfg_trefi_wire[4] ;
wire \c0|cfg_trefi_wire[5] ;
wire \c0|cfg_trefi_wire[6] ;
wire \c0|cfg_trefi_wire[7] ;
wire \c0|cfg_trefi_wire[8] ;
wire \c0|cfg_trefi_wire[9] ;
wire \c0|cfg_trefi_wire[10] ;
wire \c0|cfg_trefi_wire[11] ;
wire \c0|cfg_trefi_wire[12] ;
wire \c0|cfg_trfc_wire[0] ;
wire \c0|cfg_trfc_wire[1] ;
wire \c0|cfg_trfc_wire[2] ;
wire \c0|cfg_trfc_wire[3] ;
wire \c0|cfg_trfc_wire[4] ;
wire \c0|cfg_trfc_wire[5] ;
wire \c0|cfg_trfc_wire[6] ;
wire \c0|cfg_trfc_wire[7] ;
wire \c0|cfg_twr_wire[0] ;
wire \c0|cfg_twr_wire[1] ;
wire \c0|cfg_twr_wire[2] ;
wire \c0|cfg_twr_wire[3] ;
wire \c0|afi_mem_clk_disable[0] ;
wire \c0|cfg_dramconfig_wire[0] ;
wire \c0|cfg_dramconfig_wire[1] ;
wire \c0|cfg_dramconfig_wire[2] ;
wire \c0|cfg_dramconfig_wire[3] ;
wire \c0|cfg_dramconfig_wire[4] ;
wire \c0|cfg_dramconfig_wire[5] ;
wire \c0|cfg_dramconfig_wire[6] ;
wire \c0|cfg_dramconfig_wire[7] ;
wire \c0|cfg_dramconfig_wire[8] ;
wire \c0|cfg_dramconfig_wire[9] ;
wire \c0|cfg_dramconfig_wire[10] ;
wire \c0|cfg_dramconfig_wire[11] ;
wire \c0|cfg_dramconfig_wire[12] ;
wire \c0|cfg_dramconfig_wire[13] ;
wire \c0|cfg_dramconfig_wire[14] ;
wire \c0|cfg_dramconfig_wire[15] ;
wire \c0|cfg_dramconfig_wire[16] ;
wire \c0|cfg_dramconfig_wire[17] ;
wire \c0|cfg_dramconfig_wire[18] ;
wire \c0|cfg_dramconfig_wire[19] ;
wire \c0|cfg_dramconfig_wire[20] ;
wire \p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ;
wire \dll|dll_delayctrl[0] ;
wire \dll|dll_delayctrl[1] ;
wire \dll|dll_delayctrl[2] ;
wire \dll|dll_delayctrl[3] ;
wire \dll|dll_delayctrl[4] ;
wire \dll|dll_delayctrl[5] ;
wire \dll|dll_delayctrl[6] ;


system_altera_mem_if_oct_cyclonev oct(
	.parallelterminationcontrol({parallelterminationcontrol_15,parallelterminationcontrol_14,parallelterminationcontrol_13,parallelterminationcontrol_12,parallelterminationcontrol_11,parallelterminationcontrol_10,parallelterminationcontrol_9,parallelterminationcontrol_8,
parallelterminationcontrol_7,parallelterminationcontrol_6,parallelterminationcontrol_5,parallelterminationcontrol_4,parallelterminationcontrol_3,parallelterminationcontrol_2,parallelterminationcontrol_1,parallelterminationcontrol_0}),
	.seriesterminationcontrol({seriesterminationcontrol_15,seriesterminationcontrol_14,seriesterminationcontrol_13,seriesterminationcontrol_12,seriesterminationcontrol_11,seriesterminationcontrol_10,seriesterminationcontrol_9,seriesterminationcontrol_8,seriesterminationcontrol_7,
seriesterminationcontrol_6,seriesterminationcontrol_5,seriesterminationcontrol_4,seriesterminationcontrol_3,seriesterminationcontrol_2,seriesterminationcontrol_1,seriesterminationcontrol_0}),
	.oct_rzqin(memory_oct_rzqin));

system_altera_mem_if_dll_cyclonev dll(
	.clk(\pll|pll_write_clk ),
	.dll_delayctrl({\dll|dll_delayctrl[6] ,\dll|dll_delayctrl[5] ,\dll|dll_delayctrl[4] ,\dll|dll_delayctrl[3] ,\dll|dll_delayctrl[2] ,\dll|dll_delayctrl[1] ,\dll|dll_delayctrl[0] }));

system_altera_mem_if_hard_memory_controller_top_cyclonev c0(
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid({\p0|umemphy|afi_rdata_valid[0] }),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata({\p0|umemphy|afi_rdata[79] ,\p0|umemphy|afi_rdata[78] ,\p0|umemphy|afi_rdata[77] ,\p0|umemphy|afi_rdata[76] ,\p0|umemphy|afi_rdata[75] ,\p0|umemphy|afi_rdata[74] ,\p0|umemphy|afi_rdata[73] ,\p0|umemphy|afi_rdata[72] ,\p0|umemphy|afi_rdata[71] ,
\p0|umemphy|afi_rdata[70] ,\p0|umemphy|afi_rdata[69] ,\p0|umemphy|afi_rdata[68] ,\p0|umemphy|afi_rdata[67] ,\p0|umemphy|afi_rdata[66] ,\p0|umemphy|afi_rdata[65] ,\p0|umemphy|afi_rdata[64] ,\p0|umemphy|afi_rdata[63] ,\p0|umemphy|afi_rdata[62] ,
\p0|umemphy|afi_rdata[61] ,\p0|umemphy|afi_rdata[60] ,\p0|umemphy|afi_rdata[59] ,\p0|umemphy|afi_rdata[58] ,\p0|umemphy|afi_rdata[57] ,\p0|umemphy|afi_rdata[56] ,\p0|umemphy|afi_rdata[55] ,\p0|umemphy|afi_rdata[54] ,\p0|umemphy|afi_rdata[53] ,
\p0|umemphy|afi_rdata[52] ,\p0|umemphy|afi_rdata[51] ,\p0|umemphy|afi_rdata[50] ,\p0|umemphy|afi_rdata[49] ,\p0|umemphy|afi_rdata[48] ,\p0|umemphy|afi_rdata[47] ,\p0|umemphy|afi_rdata[46] ,\p0|umemphy|afi_rdata[45] ,\p0|umemphy|afi_rdata[44] ,
\p0|umemphy|afi_rdata[43] ,\p0|umemphy|afi_rdata[42] ,\p0|umemphy|afi_rdata[41] ,\p0|umemphy|afi_rdata[40] ,\p0|umemphy|afi_rdata[39] ,\p0|umemphy|afi_rdata[38] ,\p0|umemphy|afi_rdata[37] ,\p0|umemphy|afi_rdata[36] ,\p0|umemphy|afi_rdata[35] ,
\p0|umemphy|afi_rdata[34] ,\p0|umemphy|afi_rdata[33] ,\p0|umemphy|afi_rdata[32] ,\p0|umemphy|afi_rdata[31] ,\p0|umemphy|afi_rdata[30] ,\p0|umemphy|afi_rdata[29] ,\p0|umemphy|afi_rdata[28] ,\p0|umemphy|afi_rdata[27] ,\p0|umemphy|afi_rdata[26] ,
\p0|umemphy|afi_rdata[25] ,\p0|umemphy|afi_rdata[24] ,\p0|umemphy|afi_rdata[23] ,\p0|umemphy|afi_rdata[22] ,\p0|umemphy|afi_rdata[21] ,\p0|umemphy|afi_rdata[20] ,\p0|umemphy|afi_rdata[19] ,\p0|umemphy|afi_rdata[18] ,\p0|umemphy|afi_rdata[17] ,
\p0|umemphy|afi_rdata[16] ,\p0|umemphy|afi_rdata[15] ,\p0|umemphy|afi_rdata[14] ,\p0|umemphy|afi_rdata[13] ,\p0|umemphy|afi_rdata[12] ,\p0|umemphy|afi_rdata[11] ,\p0|umemphy|afi_rdata[10] ,\p0|umemphy|afi_rdata[9] ,\p0|umemphy|afi_rdata[8] ,
\p0|umemphy|afi_rdata[7] ,\p0|umemphy|afi_rdata[6] ,\p0|umemphy|afi_rdata[5] ,\p0|umemphy|afi_rdata[4] ,\p0|umemphy|afi_rdata[3] ,\p0|umemphy|afi_rdata[2] ,\p0|umemphy|afi_rdata[1] ,\p0|umemphy|afi_rdata[0] }),
	.afi_wlat({\p0|umemphy|afi_wlat[3] ,\p0|umemphy|afi_wlat[2] ,\p0|umemphy|afi_wlat[1] ,\p0|umemphy|afi_wlat[0] }),
	.afi_cas_n({\c0|afi_cas_n[0] }),
	.afi_ras_n({\c0|afi_ras_n[0] }),
	.afi_rst_n({\c0|afi_rst_n[0] }),
	.afi_we_n({\c0|afi_we_n[0] }),
	.afi_addr({\c0|afi_addr[19] ,\c0|afi_addr[18] ,\c0|afi_addr[17] ,\c0|afi_addr[16] ,\c0|afi_addr[15] ,\c0|afi_addr[14] ,\c0|afi_addr[13] ,\c0|afi_addr[12] ,\c0|afi_addr[11] ,\c0|afi_addr[10] ,\c0|afi_addr[9] ,\c0|afi_addr[8] ,\c0|afi_addr[7] ,\c0|afi_addr[6] ,\c0|afi_addr[5] ,
\c0|afi_addr[4] ,\c0|afi_addr[3] ,\c0|afi_addr[2] ,\c0|afi_addr[1] ,\c0|afi_addr[0] }),
	.afi_ba({\c0|afi_ba[2] ,\c0|afi_ba[1] ,\c0|afi_ba[0] }),
	.afi_cke({\c0|afi_cke[1] ,\c0|afi_cke[0] }),
	.afi_cs_n({\c0|afi_cs_n[1] ,\c0|afi_cs_n[0] }),
	.afi_dm({\c0|afi_dm_int[9] ,\c0|afi_dm_int[8] ,\c0|afi_dm_int[7] ,\c0|afi_dm_int[6] ,\c0|afi_dm_int[5] ,\c0|afi_dm_int[4] ,\c0|afi_dm_int[3] ,\c0|afi_dm_int[2] ,\c0|afi_dm_int[1] ,\c0|afi_dm_int[0] }),
	.afi_dqs_burst({\c0|afi_dqs_burst[4] ,\c0|afi_dqs_burst[3] ,\c0|afi_dqs_burst[2] ,\c0|afi_dqs_burst[1] ,\c0|afi_dqs_burst[0] }),
	.afi_odt({\c0|afi_odt[1] ,\c0|afi_odt[0] }),
	.afi_rdata_en({\c0|afi_rdata_en[4] ,\c0|afi_rdata_en[3] ,\c0|afi_rdata_en[2] ,\c0|afi_rdata_en[1] ,\c0|afi_rdata_en[0] }),
	.afi_rdata_en_full({\c0|afi_rdata_en_full[4] ,\c0|afi_rdata_en_full[3] ,\c0|afi_rdata_en_full[2] ,\c0|afi_rdata_en_full[1] ,\c0|afi_rdata_en_full[0] }),
	.afi_wdata({\c0|afi_wdata_int[79] ,\c0|afi_wdata_int[78] ,\c0|afi_wdata_int[77] ,\c0|afi_wdata_int[76] ,\c0|afi_wdata_int[75] ,\c0|afi_wdata_int[74] ,\c0|afi_wdata_int[73] ,\c0|afi_wdata_int[72] ,\c0|afi_wdata_int[71] ,\c0|afi_wdata_int[70] ,\c0|afi_wdata_int[69] ,
\c0|afi_wdata_int[68] ,\c0|afi_wdata_int[67] ,\c0|afi_wdata_int[66] ,\c0|afi_wdata_int[65] ,\c0|afi_wdata_int[64] ,\c0|afi_wdata_int[63] ,\c0|afi_wdata_int[62] ,\c0|afi_wdata_int[61] ,\c0|afi_wdata_int[60] ,\c0|afi_wdata_int[59] ,\c0|afi_wdata_int[58] ,
\c0|afi_wdata_int[57] ,\c0|afi_wdata_int[56] ,\c0|afi_wdata_int[55] ,\c0|afi_wdata_int[54] ,\c0|afi_wdata_int[53] ,\c0|afi_wdata_int[52] ,\c0|afi_wdata_int[51] ,\c0|afi_wdata_int[50] ,\c0|afi_wdata_int[49] ,\c0|afi_wdata_int[48] ,\c0|afi_wdata_int[47] ,
\c0|afi_wdata_int[46] ,\c0|afi_wdata_int[45] ,\c0|afi_wdata_int[44] ,\c0|afi_wdata_int[43] ,\c0|afi_wdata_int[42] ,\c0|afi_wdata_int[41] ,\c0|afi_wdata_int[40] ,\c0|afi_wdata_int[39] ,\c0|afi_wdata_int[38] ,\c0|afi_wdata_int[37] ,\c0|afi_wdata_int[36] ,
\c0|afi_wdata_int[35] ,\c0|afi_wdata_int[34] ,\c0|afi_wdata_int[33] ,\c0|afi_wdata_int[32] ,\c0|afi_wdata_int[31] ,\c0|afi_wdata_int[30] ,\c0|afi_wdata_int[29] ,\c0|afi_wdata_int[28] ,\c0|afi_wdata_int[27] ,\c0|afi_wdata_int[26] ,\c0|afi_wdata_int[25] ,
\c0|afi_wdata_int[24] ,\c0|afi_wdata_int[23] ,\c0|afi_wdata_int[22] ,\c0|afi_wdata_int[21] ,\c0|afi_wdata_int[20] ,\c0|afi_wdata_int[19] ,\c0|afi_wdata_int[18] ,\c0|afi_wdata_int[17] ,\c0|afi_wdata_int[16] ,\c0|afi_wdata_int[15] ,\c0|afi_wdata_int[14] ,
\c0|afi_wdata_int[13] ,\c0|afi_wdata_int[12] ,\c0|afi_wdata_int[11] ,\c0|afi_wdata_int[10] ,\c0|afi_wdata_int[9] ,\c0|afi_wdata_int[8] ,\c0|afi_wdata_int[7] ,\c0|afi_wdata_int[6] ,\c0|afi_wdata_int[5] ,\c0|afi_wdata_int[4] ,\c0|afi_wdata_int[3] ,\c0|afi_wdata_int[2] ,
\c0|afi_wdata_int[1] ,\c0|afi_wdata_int[0] }),
	.afi_wdata_valid({\c0|afi_wdata_valid[4] ,\c0|afi_wdata_valid[3] ,\c0|afi_wdata_valid[2] ,\c0|afi_wdata_valid[1] ,\c0|afi_wdata_valid[0] }),
	.cfg_addlat({cfg_addlat_unconnected_wire_7,cfg_addlat_unconnected_wire_6,cfg_addlat_unconnected_wire_5,\c0|cfg_addlat_wire[4] ,\c0|cfg_addlat_wire[3] ,\c0|cfg_addlat_wire[2] ,\c0|cfg_addlat_wire[1] ,\c0|cfg_addlat_wire[0] }),
	.cfg_bankaddrwidth({cfg_bankaddrwidth_unconnected_wire_7,cfg_bankaddrwidth_unconnected_wire_6,cfg_bankaddrwidth_unconnected_wire_5,cfg_bankaddrwidth_unconnected_wire_4,cfg_bankaddrwidth_unconnected_wire_3,\c0|cfg_bankaddrwidth_wire[2] ,\c0|cfg_bankaddrwidth_wire[1] ,
\c0|cfg_bankaddrwidth_wire[0] }),
	.cfg_caswrlat({cfg_caswrlat_unconnected_wire_7,cfg_caswrlat_unconnected_wire_6,cfg_caswrlat_unconnected_wire_5,cfg_caswrlat_unconnected_wire_4,\c0|cfg_caswrlat_wire[3] ,\c0|cfg_caswrlat_wire[2] ,\c0|cfg_caswrlat_wire[1] ,\c0|cfg_caswrlat_wire[0] }),
	.cfg_coladdrwidth({cfg_coladdrwidth_unconnected_wire_7,cfg_coladdrwidth_unconnected_wire_6,cfg_coladdrwidth_unconnected_wire_5,\c0|cfg_coladdrwidth_wire[4] ,\c0|cfg_coladdrwidth_wire[3] ,\c0|cfg_coladdrwidth_wire[2] ,\c0|cfg_coladdrwidth_wire[1] ,\c0|cfg_coladdrwidth_wire[0] }),
	.cfg_csaddrwidth({cfg_csaddrwidth_unconnected_wire_7,cfg_csaddrwidth_unconnected_wire_6,cfg_csaddrwidth_unconnected_wire_5,cfg_csaddrwidth_unconnected_wire_4,cfg_csaddrwidth_unconnected_wire_3,\c0|cfg_csaddrwidth_wire[2] ,\c0|cfg_csaddrwidth_wire[1] ,\c0|cfg_csaddrwidth_wire[0] }),
	.cfg_devicewidth({cfg_devicewidth_unconnected_wire_7,cfg_devicewidth_unconnected_wire_6,cfg_devicewidth_unconnected_wire_5,cfg_devicewidth_unconnected_wire_4,\c0|cfg_devicewidth_wire[3] ,\c0|cfg_devicewidth_wire[2] ,\c0|cfg_devicewidth_wire[1] ,\c0|cfg_devicewidth_wire[0] }),
	.cfg_interfacewidth({\c0|cfg_interfacewidth_wire[7] ,\c0|cfg_interfacewidth_wire[6] ,\c0|cfg_interfacewidth_wire[5] ,\c0|cfg_interfacewidth_wire[4] ,\c0|cfg_interfacewidth_wire[3] ,\c0|cfg_interfacewidth_wire[2] ,\c0|cfg_interfacewidth_wire[1] ,\c0|cfg_interfacewidth_wire[0] }),
	.cfg_rowaddrwidth({cfg_rowaddrwidth_unconnected_wire_7,cfg_rowaddrwidth_unconnected_wire_6,cfg_rowaddrwidth_unconnected_wire_5,\c0|cfg_rowaddrwidth_wire[4] ,\c0|cfg_rowaddrwidth_wire[3] ,\c0|cfg_rowaddrwidth_wire[2] ,\c0|cfg_rowaddrwidth_wire[1] ,\c0|cfg_rowaddrwidth_wire[0] }),
	.cfg_tcl({cfg_tcl_unconnected_wire_7,cfg_tcl_unconnected_wire_6,cfg_tcl_unconnected_wire_5,\c0|cfg_tcl_wire[4] ,\c0|cfg_tcl_wire[3] ,\c0|cfg_tcl_wire[2] ,\c0|cfg_tcl_wire[1] ,\c0|cfg_tcl_wire[0] }),
	.cfg_tmrd({cfg_tmrd_unconnected_wire_7,cfg_tmrd_unconnected_wire_6,cfg_tmrd_unconnected_wire_5,cfg_tmrd_unconnected_wire_4,\c0|cfg_tmrd_wire[3] ,\c0|cfg_tmrd_wire[2] ,\c0|cfg_tmrd_wire[1] ,\c0|cfg_tmrd_wire[0] }),
	.cfg_trefi({cfg_trefi_unconnected_wire_15,cfg_trefi_unconnected_wire_14,cfg_trefi_unconnected_wire_13,\c0|cfg_trefi_wire[12] ,\c0|cfg_trefi_wire[11] ,\c0|cfg_trefi_wire[10] ,\c0|cfg_trefi_wire[9] ,\c0|cfg_trefi_wire[8] ,\c0|cfg_trefi_wire[7] ,\c0|cfg_trefi_wire[6] ,
\c0|cfg_trefi_wire[5] ,\c0|cfg_trefi_wire[4] ,\c0|cfg_trefi_wire[3] ,\c0|cfg_trefi_wire[2] ,\c0|cfg_trefi_wire[1] ,\c0|cfg_trefi_wire[0] }),
	.cfg_trfc({\c0|cfg_trfc_wire[7] ,\c0|cfg_trfc_wire[6] ,\c0|cfg_trfc_wire[5] ,\c0|cfg_trfc_wire[4] ,\c0|cfg_trfc_wire[3] ,\c0|cfg_trfc_wire[2] ,\c0|cfg_trfc_wire[1] ,\c0|cfg_trfc_wire[0] }),
	.cfg_twr({cfg_twr_unconnected_wire_7,cfg_twr_unconnected_wire_6,cfg_twr_unconnected_wire_5,cfg_twr_unconnected_wire_4,\c0|cfg_twr_wire[3] ,\c0|cfg_twr_wire[2] ,\c0|cfg_twr_wire[1] ,\c0|cfg_twr_wire[0] }),
	.afi_mem_clk_disable({\c0|afi_mem_clk_disable[0] }),
	.cfg_dramconfig({cfg_dramconfig_unconnected_wire_23,cfg_dramconfig_unconnected_wire_22,cfg_dramconfig_unconnected_wire_21,\c0|cfg_dramconfig_wire[20] ,\c0|cfg_dramconfig_wire[19] ,\c0|cfg_dramconfig_wire[18] ,\c0|cfg_dramconfig_wire[17] ,\c0|cfg_dramconfig_wire[16] ,
\c0|cfg_dramconfig_wire[15] ,\c0|cfg_dramconfig_wire[14] ,\c0|cfg_dramconfig_wire[13] ,\c0|cfg_dramconfig_wire[12] ,\c0|cfg_dramconfig_wire[11] ,\c0|cfg_dramconfig_wire[10] ,\c0|cfg_dramconfig_wire[9] ,\c0|cfg_dramconfig_wire[8] ,\c0|cfg_dramconfig_wire[7] ,
\c0|cfg_dramconfig_wire[6] ,\c0|cfg_dramconfig_wire[5] ,\c0|cfg_dramconfig_wire[4] ,\c0|cfg_dramconfig_wire[3] ,\c0|cfg_dramconfig_wire[2] ,\c0|cfg_dramconfig_wire[1] ,\c0|cfg_dramconfig_wire[0] }),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ));

system_hps_sdram_p0 p0(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid_0(\p0|umemphy|afi_rdata_valid[0] ),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata_0(\p0|umemphy|afi_rdata[0] ),
	.afi_rdata_1(\p0|umemphy|afi_rdata[1] ),
	.afi_rdata_2(\p0|umemphy|afi_rdata[2] ),
	.afi_rdata_3(\p0|umemphy|afi_rdata[3] ),
	.afi_rdata_4(\p0|umemphy|afi_rdata[4] ),
	.afi_rdata_5(\p0|umemphy|afi_rdata[5] ),
	.afi_rdata_6(\p0|umemphy|afi_rdata[6] ),
	.afi_rdata_7(\p0|umemphy|afi_rdata[7] ),
	.afi_rdata_8(\p0|umemphy|afi_rdata[8] ),
	.afi_rdata_9(\p0|umemphy|afi_rdata[9] ),
	.afi_rdata_10(\p0|umemphy|afi_rdata[10] ),
	.afi_rdata_11(\p0|umemphy|afi_rdata[11] ),
	.afi_rdata_12(\p0|umemphy|afi_rdata[12] ),
	.afi_rdata_13(\p0|umemphy|afi_rdata[13] ),
	.afi_rdata_14(\p0|umemphy|afi_rdata[14] ),
	.afi_rdata_15(\p0|umemphy|afi_rdata[15] ),
	.afi_rdata_16(\p0|umemphy|afi_rdata[16] ),
	.afi_rdata_17(\p0|umemphy|afi_rdata[17] ),
	.afi_rdata_18(\p0|umemphy|afi_rdata[18] ),
	.afi_rdata_19(\p0|umemphy|afi_rdata[19] ),
	.afi_rdata_20(\p0|umemphy|afi_rdata[20] ),
	.afi_rdata_21(\p0|umemphy|afi_rdata[21] ),
	.afi_rdata_22(\p0|umemphy|afi_rdata[22] ),
	.afi_rdata_23(\p0|umemphy|afi_rdata[23] ),
	.afi_rdata_24(\p0|umemphy|afi_rdata[24] ),
	.afi_rdata_25(\p0|umemphy|afi_rdata[25] ),
	.afi_rdata_26(\p0|umemphy|afi_rdata[26] ),
	.afi_rdata_27(\p0|umemphy|afi_rdata[27] ),
	.afi_rdata_28(\p0|umemphy|afi_rdata[28] ),
	.afi_rdata_29(\p0|umemphy|afi_rdata[29] ),
	.afi_rdata_30(\p0|umemphy|afi_rdata[30] ),
	.afi_rdata_31(\p0|umemphy|afi_rdata[31] ),
	.afi_rdata_32(\p0|umemphy|afi_rdata[32] ),
	.afi_rdata_33(\p0|umemphy|afi_rdata[33] ),
	.afi_rdata_34(\p0|umemphy|afi_rdata[34] ),
	.afi_rdata_35(\p0|umemphy|afi_rdata[35] ),
	.afi_rdata_36(\p0|umemphy|afi_rdata[36] ),
	.afi_rdata_37(\p0|umemphy|afi_rdata[37] ),
	.afi_rdata_38(\p0|umemphy|afi_rdata[38] ),
	.afi_rdata_39(\p0|umemphy|afi_rdata[39] ),
	.afi_rdata_40(\p0|umemphy|afi_rdata[40] ),
	.afi_rdata_41(\p0|umemphy|afi_rdata[41] ),
	.afi_rdata_42(\p0|umemphy|afi_rdata[42] ),
	.afi_rdata_43(\p0|umemphy|afi_rdata[43] ),
	.afi_rdata_44(\p0|umemphy|afi_rdata[44] ),
	.afi_rdata_45(\p0|umemphy|afi_rdata[45] ),
	.afi_rdata_46(\p0|umemphy|afi_rdata[46] ),
	.afi_rdata_47(\p0|umemphy|afi_rdata[47] ),
	.afi_rdata_48(\p0|umemphy|afi_rdata[48] ),
	.afi_rdata_49(\p0|umemphy|afi_rdata[49] ),
	.afi_rdata_50(\p0|umemphy|afi_rdata[50] ),
	.afi_rdata_51(\p0|umemphy|afi_rdata[51] ),
	.afi_rdata_52(\p0|umemphy|afi_rdata[52] ),
	.afi_rdata_53(\p0|umemphy|afi_rdata[53] ),
	.afi_rdata_54(\p0|umemphy|afi_rdata[54] ),
	.afi_rdata_55(\p0|umemphy|afi_rdata[55] ),
	.afi_rdata_56(\p0|umemphy|afi_rdata[56] ),
	.afi_rdata_57(\p0|umemphy|afi_rdata[57] ),
	.afi_rdata_58(\p0|umemphy|afi_rdata[58] ),
	.afi_rdata_59(\p0|umemphy|afi_rdata[59] ),
	.afi_rdata_60(\p0|umemphy|afi_rdata[60] ),
	.afi_rdata_61(\p0|umemphy|afi_rdata[61] ),
	.afi_rdata_62(\p0|umemphy|afi_rdata[62] ),
	.afi_rdata_63(\p0|umemphy|afi_rdata[63] ),
	.afi_rdata_64(\p0|umemphy|afi_rdata[64] ),
	.afi_rdata_65(\p0|umemphy|afi_rdata[65] ),
	.afi_rdata_66(\p0|umemphy|afi_rdata[66] ),
	.afi_rdata_67(\p0|umemphy|afi_rdata[67] ),
	.afi_rdata_68(\p0|umemphy|afi_rdata[68] ),
	.afi_rdata_69(\p0|umemphy|afi_rdata[69] ),
	.afi_rdata_70(\p0|umemphy|afi_rdata[70] ),
	.afi_rdata_71(\p0|umemphy|afi_rdata[71] ),
	.afi_rdata_72(\p0|umemphy|afi_rdata[72] ),
	.afi_rdata_73(\p0|umemphy|afi_rdata[73] ),
	.afi_rdata_74(\p0|umemphy|afi_rdata[74] ),
	.afi_rdata_75(\p0|umemphy|afi_rdata[75] ),
	.afi_rdata_76(\p0|umemphy|afi_rdata[76] ),
	.afi_rdata_77(\p0|umemphy|afi_rdata[77] ),
	.afi_rdata_78(\p0|umemphy|afi_rdata[78] ),
	.afi_rdata_79(\p0|umemphy|afi_rdata[79] ),
	.afi_wlat_0(\p0|umemphy|afi_wlat[0] ),
	.afi_wlat_1(\p0|umemphy|afi_wlat[1] ),
	.afi_wlat_2(\p0|umemphy|afi_wlat[2] ),
	.afi_wlat_3(\p0|umemphy|afi_wlat[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n_0(\c0|afi_cas_n[0] ),
	.afi_ras_n_0(\c0|afi_ras_n[0] ),
	.afi_rst_n_0(\c0|afi_rst_n[0] ),
	.afi_we_n_0(\c0|afi_we_n[0] ),
	.afi_addr_0(\c0|afi_addr[0] ),
	.afi_addr_1(\c0|afi_addr[1] ),
	.afi_addr_2(\c0|afi_addr[2] ),
	.afi_addr_3(\c0|afi_addr[3] ),
	.afi_addr_4(\c0|afi_addr[4] ),
	.afi_addr_5(\c0|afi_addr[5] ),
	.afi_addr_6(\c0|afi_addr[6] ),
	.afi_addr_7(\c0|afi_addr[7] ),
	.afi_addr_8(\c0|afi_addr[8] ),
	.afi_addr_9(\c0|afi_addr[9] ),
	.afi_addr_10(\c0|afi_addr[10] ),
	.afi_addr_11(\c0|afi_addr[11] ),
	.afi_addr_12(\c0|afi_addr[12] ),
	.afi_addr_13(\c0|afi_addr[13] ),
	.afi_addr_14(\c0|afi_addr[14] ),
	.afi_addr_15(\c0|afi_addr[15] ),
	.afi_addr_16(\c0|afi_addr[16] ),
	.afi_addr_17(\c0|afi_addr[17] ),
	.afi_addr_18(\c0|afi_addr[18] ),
	.afi_addr_19(\c0|afi_addr[19] ),
	.afi_ba_0(\c0|afi_ba[0] ),
	.afi_ba_1(\c0|afi_ba[1] ),
	.afi_ba_2(\c0|afi_ba[2] ),
	.afi_cke_0(\c0|afi_cke[0] ),
	.afi_cke_1(\c0|afi_cke[1] ),
	.afi_cs_n_0(\c0|afi_cs_n[0] ),
	.afi_cs_n_1(\c0|afi_cs_n[1] ),
	.afi_dm_int_0(\c0|afi_dm_int[0] ),
	.afi_dm_int_1(\c0|afi_dm_int[1] ),
	.afi_dm_int_2(\c0|afi_dm_int[2] ),
	.afi_dm_int_3(\c0|afi_dm_int[3] ),
	.afi_dm_int_4(\c0|afi_dm_int[4] ),
	.afi_dm_int_5(\c0|afi_dm_int[5] ),
	.afi_dm_int_6(\c0|afi_dm_int[6] ),
	.afi_dm_int_7(\c0|afi_dm_int[7] ),
	.afi_dm_int_8(\c0|afi_dm_int[8] ),
	.afi_dm_int_9(\c0|afi_dm_int[9] ),
	.afi_dqs_burst_0(\c0|afi_dqs_burst[0] ),
	.afi_dqs_burst_1(\c0|afi_dqs_burst[1] ),
	.afi_dqs_burst_2(\c0|afi_dqs_burst[2] ),
	.afi_dqs_burst_3(\c0|afi_dqs_burst[3] ),
	.afi_dqs_burst_4(\c0|afi_dqs_burst[4] ),
	.afi_odt_0(\c0|afi_odt[0] ),
	.afi_odt_1(\c0|afi_odt[1] ),
	.afi_rdata_en_0(\c0|afi_rdata_en[0] ),
	.afi_rdata_en_1(\c0|afi_rdata_en[1] ),
	.afi_rdata_en_2(\c0|afi_rdata_en[2] ),
	.afi_rdata_en_3(\c0|afi_rdata_en[3] ),
	.afi_rdata_en_4(\c0|afi_rdata_en[4] ),
	.afi_rdata_en_full_0(\c0|afi_rdata_en_full[0] ),
	.afi_rdata_en_full_1(\c0|afi_rdata_en_full[1] ),
	.afi_rdata_en_full_2(\c0|afi_rdata_en_full[2] ),
	.afi_rdata_en_full_3(\c0|afi_rdata_en_full[3] ),
	.afi_rdata_en_full_4(\c0|afi_rdata_en_full[4] ),
	.afi_wdata_int_0(\c0|afi_wdata_int[0] ),
	.afi_wdata_int_1(\c0|afi_wdata_int[1] ),
	.afi_wdata_int_2(\c0|afi_wdata_int[2] ),
	.afi_wdata_int_3(\c0|afi_wdata_int[3] ),
	.afi_wdata_int_4(\c0|afi_wdata_int[4] ),
	.afi_wdata_int_5(\c0|afi_wdata_int[5] ),
	.afi_wdata_int_6(\c0|afi_wdata_int[6] ),
	.afi_wdata_int_7(\c0|afi_wdata_int[7] ),
	.afi_wdata_int_8(\c0|afi_wdata_int[8] ),
	.afi_wdata_int_9(\c0|afi_wdata_int[9] ),
	.afi_wdata_int_10(\c0|afi_wdata_int[10] ),
	.afi_wdata_int_11(\c0|afi_wdata_int[11] ),
	.afi_wdata_int_12(\c0|afi_wdata_int[12] ),
	.afi_wdata_int_13(\c0|afi_wdata_int[13] ),
	.afi_wdata_int_14(\c0|afi_wdata_int[14] ),
	.afi_wdata_int_15(\c0|afi_wdata_int[15] ),
	.afi_wdata_int_16(\c0|afi_wdata_int[16] ),
	.afi_wdata_int_17(\c0|afi_wdata_int[17] ),
	.afi_wdata_int_18(\c0|afi_wdata_int[18] ),
	.afi_wdata_int_19(\c0|afi_wdata_int[19] ),
	.afi_wdata_int_20(\c0|afi_wdata_int[20] ),
	.afi_wdata_int_21(\c0|afi_wdata_int[21] ),
	.afi_wdata_int_22(\c0|afi_wdata_int[22] ),
	.afi_wdata_int_23(\c0|afi_wdata_int[23] ),
	.afi_wdata_int_24(\c0|afi_wdata_int[24] ),
	.afi_wdata_int_25(\c0|afi_wdata_int[25] ),
	.afi_wdata_int_26(\c0|afi_wdata_int[26] ),
	.afi_wdata_int_27(\c0|afi_wdata_int[27] ),
	.afi_wdata_int_28(\c0|afi_wdata_int[28] ),
	.afi_wdata_int_29(\c0|afi_wdata_int[29] ),
	.afi_wdata_int_30(\c0|afi_wdata_int[30] ),
	.afi_wdata_int_31(\c0|afi_wdata_int[31] ),
	.afi_wdata_int_32(\c0|afi_wdata_int[32] ),
	.afi_wdata_int_33(\c0|afi_wdata_int[33] ),
	.afi_wdata_int_34(\c0|afi_wdata_int[34] ),
	.afi_wdata_int_35(\c0|afi_wdata_int[35] ),
	.afi_wdata_int_36(\c0|afi_wdata_int[36] ),
	.afi_wdata_int_37(\c0|afi_wdata_int[37] ),
	.afi_wdata_int_38(\c0|afi_wdata_int[38] ),
	.afi_wdata_int_39(\c0|afi_wdata_int[39] ),
	.afi_wdata_int_40(\c0|afi_wdata_int[40] ),
	.afi_wdata_int_41(\c0|afi_wdata_int[41] ),
	.afi_wdata_int_42(\c0|afi_wdata_int[42] ),
	.afi_wdata_int_43(\c0|afi_wdata_int[43] ),
	.afi_wdata_int_44(\c0|afi_wdata_int[44] ),
	.afi_wdata_int_45(\c0|afi_wdata_int[45] ),
	.afi_wdata_int_46(\c0|afi_wdata_int[46] ),
	.afi_wdata_int_47(\c0|afi_wdata_int[47] ),
	.afi_wdata_int_48(\c0|afi_wdata_int[48] ),
	.afi_wdata_int_49(\c0|afi_wdata_int[49] ),
	.afi_wdata_int_50(\c0|afi_wdata_int[50] ),
	.afi_wdata_int_51(\c0|afi_wdata_int[51] ),
	.afi_wdata_int_52(\c0|afi_wdata_int[52] ),
	.afi_wdata_int_53(\c0|afi_wdata_int[53] ),
	.afi_wdata_int_54(\c0|afi_wdata_int[54] ),
	.afi_wdata_int_55(\c0|afi_wdata_int[55] ),
	.afi_wdata_int_56(\c0|afi_wdata_int[56] ),
	.afi_wdata_int_57(\c0|afi_wdata_int[57] ),
	.afi_wdata_int_58(\c0|afi_wdata_int[58] ),
	.afi_wdata_int_59(\c0|afi_wdata_int[59] ),
	.afi_wdata_int_60(\c0|afi_wdata_int[60] ),
	.afi_wdata_int_61(\c0|afi_wdata_int[61] ),
	.afi_wdata_int_62(\c0|afi_wdata_int[62] ),
	.afi_wdata_int_63(\c0|afi_wdata_int[63] ),
	.afi_wdata_int_64(\c0|afi_wdata_int[64] ),
	.afi_wdata_int_65(\c0|afi_wdata_int[65] ),
	.afi_wdata_int_66(\c0|afi_wdata_int[66] ),
	.afi_wdata_int_67(\c0|afi_wdata_int[67] ),
	.afi_wdata_int_68(\c0|afi_wdata_int[68] ),
	.afi_wdata_int_69(\c0|afi_wdata_int[69] ),
	.afi_wdata_int_70(\c0|afi_wdata_int[70] ),
	.afi_wdata_int_71(\c0|afi_wdata_int[71] ),
	.afi_wdata_int_72(\c0|afi_wdata_int[72] ),
	.afi_wdata_int_73(\c0|afi_wdata_int[73] ),
	.afi_wdata_int_74(\c0|afi_wdata_int[74] ),
	.afi_wdata_int_75(\c0|afi_wdata_int[75] ),
	.afi_wdata_int_76(\c0|afi_wdata_int[76] ),
	.afi_wdata_int_77(\c0|afi_wdata_int[77] ),
	.afi_wdata_int_78(\c0|afi_wdata_int[78] ),
	.afi_wdata_int_79(\c0|afi_wdata_int[79] ),
	.afi_wdata_valid_0(\c0|afi_wdata_valid[0] ),
	.afi_wdata_valid_1(\c0|afi_wdata_valid[1] ),
	.afi_wdata_valid_2(\c0|afi_wdata_valid[2] ),
	.afi_wdata_valid_3(\c0|afi_wdata_valid[3] ),
	.afi_wdata_valid_4(\c0|afi_wdata_valid[4] ),
	.cfg_addlat_wire_0(\c0|cfg_addlat_wire[0] ),
	.cfg_addlat_wire_1(\c0|cfg_addlat_wire[1] ),
	.cfg_addlat_wire_2(\c0|cfg_addlat_wire[2] ),
	.cfg_addlat_wire_3(\c0|cfg_addlat_wire[3] ),
	.cfg_addlat_wire_4(\c0|cfg_addlat_wire[4] ),
	.cfg_bankaddrwidth_wire_0(\c0|cfg_bankaddrwidth_wire[0] ),
	.cfg_bankaddrwidth_wire_1(\c0|cfg_bankaddrwidth_wire[1] ),
	.cfg_bankaddrwidth_wire_2(\c0|cfg_bankaddrwidth_wire[2] ),
	.cfg_caswrlat_wire_0(\c0|cfg_caswrlat_wire[0] ),
	.cfg_caswrlat_wire_1(\c0|cfg_caswrlat_wire[1] ),
	.cfg_caswrlat_wire_2(\c0|cfg_caswrlat_wire[2] ),
	.cfg_caswrlat_wire_3(\c0|cfg_caswrlat_wire[3] ),
	.cfg_coladdrwidth_wire_0(\c0|cfg_coladdrwidth_wire[0] ),
	.cfg_coladdrwidth_wire_1(\c0|cfg_coladdrwidth_wire[1] ),
	.cfg_coladdrwidth_wire_2(\c0|cfg_coladdrwidth_wire[2] ),
	.cfg_coladdrwidth_wire_3(\c0|cfg_coladdrwidth_wire[3] ),
	.cfg_coladdrwidth_wire_4(\c0|cfg_coladdrwidth_wire[4] ),
	.cfg_csaddrwidth_wire_0(\c0|cfg_csaddrwidth_wire[0] ),
	.cfg_csaddrwidth_wire_1(\c0|cfg_csaddrwidth_wire[1] ),
	.cfg_csaddrwidth_wire_2(\c0|cfg_csaddrwidth_wire[2] ),
	.cfg_devicewidth_wire_0(\c0|cfg_devicewidth_wire[0] ),
	.cfg_devicewidth_wire_1(\c0|cfg_devicewidth_wire[1] ),
	.cfg_devicewidth_wire_2(\c0|cfg_devicewidth_wire[2] ),
	.cfg_devicewidth_wire_3(\c0|cfg_devicewidth_wire[3] ),
	.cfg_interfacewidth_wire_0(\c0|cfg_interfacewidth_wire[0] ),
	.cfg_interfacewidth_wire_1(\c0|cfg_interfacewidth_wire[1] ),
	.cfg_interfacewidth_wire_2(\c0|cfg_interfacewidth_wire[2] ),
	.cfg_interfacewidth_wire_3(\c0|cfg_interfacewidth_wire[3] ),
	.cfg_interfacewidth_wire_4(\c0|cfg_interfacewidth_wire[4] ),
	.cfg_interfacewidth_wire_5(\c0|cfg_interfacewidth_wire[5] ),
	.cfg_interfacewidth_wire_6(\c0|cfg_interfacewidth_wire[6] ),
	.cfg_interfacewidth_wire_7(\c0|cfg_interfacewidth_wire[7] ),
	.cfg_rowaddrwidth_wire_0(\c0|cfg_rowaddrwidth_wire[0] ),
	.cfg_rowaddrwidth_wire_1(\c0|cfg_rowaddrwidth_wire[1] ),
	.cfg_rowaddrwidth_wire_2(\c0|cfg_rowaddrwidth_wire[2] ),
	.cfg_rowaddrwidth_wire_3(\c0|cfg_rowaddrwidth_wire[3] ),
	.cfg_rowaddrwidth_wire_4(\c0|cfg_rowaddrwidth_wire[4] ),
	.cfg_tcl_wire_0(\c0|cfg_tcl_wire[0] ),
	.cfg_tcl_wire_1(\c0|cfg_tcl_wire[1] ),
	.cfg_tcl_wire_2(\c0|cfg_tcl_wire[2] ),
	.cfg_tcl_wire_3(\c0|cfg_tcl_wire[3] ),
	.cfg_tcl_wire_4(\c0|cfg_tcl_wire[4] ),
	.cfg_tmrd_wire_0(\c0|cfg_tmrd_wire[0] ),
	.cfg_tmrd_wire_1(\c0|cfg_tmrd_wire[1] ),
	.cfg_tmrd_wire_2(\c0|cfg_tmrd_wire[2] ),
	.cfg_tmrd_wire_3(\c0|cfg_tmrd_wire[3] ),
	.cfg_trefi_wire_0(\c0|cfg_trefi_wire[0] ),
	.cfg_trefi_wire_1(\c0|cfg_trefi_wire[1] ),
	.cfg_trefi_wire_2(\c0|cfg_trefi_wire[2] ),
	.cfg_trefi_wire_3(\c0|cfg_trefi_wire[3] ),
	.cfg_trefi_wire_4(\c0|cfg_trefi_wire[4] ),
	.cfg_trefi_wire_5(\c0|cfg_trefi_wire[5] ),
	.cfg_trefi_wire_6(\c0|cfg_trefi_wire[6] ),
	.cfg_trefi_wire_7(\c0|cfg_trefi_wire[7] ),
	.cfg_trefi_wire_8(\c0|cfg_trefi_wire[8] ),
	.cfg_trefi_wire_9(\c0|cfg_trefi_wire[9] ),
	.cfg_trefi_wire_10(\c0|cfg_trefi_wire[10] ),
	.cfg_trefi_wire_11(\c0|cfg_trefi_wire[11] ),
	.cfg_trefi_wire_12(\c0|cfg_trefi_wire[12] ),
	.cfg_trfc_wire_0(\c0|cfg_trfc_wire[0] ),
	.cfg_trfc_wire_1(\c0|cfg_trfc_wire[1] ),
	.cfg_trfc_wire_2(\c0|cfg_trfc_wire[2] ),
	.cfg_trfc_wire_3(\c0|cfg_trfc_wire[3] ),
	.cfg_trfc_wire_4(\c0|cfg_trfc_wire[4] ),
	.cfg_trfc_wire_5(\c0|cfg_trfc_wire[5] ),
	.cfg_trfc_wire_6(\c0|cfg_trfc_wire[6] ),
	.cfg_trfc_wire_7(\c0|cfg_trfc_wire[7] ),
	.cfg_twr_wire_0(\c0|cfg_twr_wire[0] ),
	.cfg_twr_wire_1(\c0|cfg_twr_wire[1] ),
	.cfg_twr_wire_2(\c0|cfg_twr_wire[2] ),
	.cfg_twr_wire_3(\c0|cfg_twr_wire[3] ),
	.afi_mem_clk_disable_0(\c0|afi_mem_clk_disable[0] ),
	.cfg_dramconfig_wire_0(\c0|cfg_dramconfig_wire[0] ),
	.cfg_dramconfig_wire_1(\c0|cfg_dramconfig_wire[1] ),
	.cfg_dramconfig_wire_2(\c0|cfg_dramconfig_wire[2] ),
	.cfg_dramconfig_wire_3(\c0|cfg_dramconfig_wire[3] ),
	.cfg_dramconfig_wire_4(\c0|cfg_dramconfig_wire[4] ),
	.cfg_dramconfig_wire_5(\c0|cfg_dramconfig_wire[5] ),
	.cfg_dramconfig_wire_6(\c0|cfg_dramconfig_wire[6] ),
	.cfg_dramconfig_wire_7(\c0|cfg_dramconfig_wire[7] ),
	.cfg_dramconfig_wire_8(\c0|cfg_dramconfig_wire[8] ),
	.cfg_dramconfig_wire_9(\c0|cfg_dramconfig_wire[9] ),
	.cfg_dramconfig_wire_10(\c0|cfg_dramconfig_wire[10] ),
	.cfg_dramconfig_wire_11(\c0|cfg_dramconfig_wire[11] ),
	.cfg_dramconfig_wire_12(\c0|cfg_dramconfig_wire[12] ),
	.cfg_dramconfig_wire_13(\c0|cfg_dramconfig_wire[13] ),
	.cfg_dramconfig_wire_14(\c0|cfg_dramconfig_wire[14] ),
	.cfg_dramconfig_wire_15(\c0|cfg_dramconfig_wire[15] ),
	.cfg_dramconfig_wire_16(\c0|cfg_dramconfig_wire[16] ),
	.cfg_dramconfig_wire_17(\c0|cfg_dramconfig_wire[17] ),
	.cfg_dramconfig_wire_18(\c0|cfg_dramconfig_wire[18] ),
	.cfg_dramconfig_wire_19(\c0|cfg_dramconfig_wire[19] ),
	.cfg_dramconfig_wire_20(\c0|cfg_dramconfig_wire[20] ),
	.leveled_dqs_clocks_0(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ),
	.dll_delayctrl_0(\dll|dll_delayctrl[0] ),
	.dll_delayctrl_1(\dll|dll_delayctrl[1] ),
	.dll_delayctrl_2(\dll|dll_delayctrl[2] ),
	.dll_delayctrl_3(\dll|dll_delayctrl[3] ),
	.dll_delayctrl_4(\dll|dll_delayctrl[4] ),
	.dll_delayctrl_5(\dll|dll_delayctrl[5] ),
	.dll_delayctrl_6(\dll|dll_delayctrl[6] ),
	.GND_port(GND_port));

system_hps_sdram_pll pll(
	.afi_half_clk(\pll|afi_clk ),
	.pll_write_clk_pre_phy_clk(\pll|pll_write_clk ));

endmodule

module system_altera_mem_if_dll_cyclonev (
	clk,
	dll_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	[6:0] dll_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [6:0] dll_wys_m_DELAYCTRLOUT_bus;

assign dll_delayctrl[0] = dll_wys_m_DELAYCTRLOUT_bus[0];
assign dll_delayctrl[1] = dll_wys_m_DELAYCTRLOUT_bus[1];
assign dll_delayctrl[2] = dll_wys_m_DELAYCTRLOUT_bus[2];
assign dll_delayctrl[3] = dll_wys_m_DELAYCTRLOUT_bus[3];
assign dll_delayctrl[4] = dll_wys_m_DELAYCTRLOUT_bus[4];
assign dll_delayctrl[5] = dll_wys_m_DELAYCTRLOUT_bus[5];
assign dll_delayctrl[6] = dll_wys_m_DELAYCTRLOUT_bus[6];

cyclonev_dll dll_wys_m(
	.clk(clk),
	.aload(vcc),
	.upndnin(gnd),
	.upndninclkena(gnd),
	.dqsupdate(),
	.upndnout(),
	.delayctrlout(dll_wys_m_DELAYCTRLOUT_bus));
defparam dll_wys_m.delayctrlout_mode = "normal";
defparam dll_wys_m.input_frequency = "2500 ps";
defparam dll_wys_m.jitter_reduction = "true";
defparam dll_wys_m.sim_buffer_delay_increment = 10;
defparam dll_wys_m.sim_buffer_intrinsic_delay = 175;
defparam dll_wys_m.sim_valid_lock = 16;
defparam dll_wys_m.sim_valid_lockcount = 0;
defparam dll_wys_m.static_delay_ctrl = 8;
defparam dll_wys_m.upndnout_mode = "clock";
defparam dll_wys_m.use_upndnin = "false";
defparam dll_wys_m.use_upndninclkena = "false";

endmodule

module system_altera_mem_if_hard_memory_controller_top_cyclonev (
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk)/* synthesis synthesis_greybox=0 */;
input 	afi_cal_fail;
input 	afi_cal_success;
input 	[0:0] afi_rdata_valid;
input 	ctl_reset_n;
input 	[79:0] afi_rdata;
input 	[3:0] afi_wlat;
output 	[0:0] afi_cas_n;
output 	[0:0] afi_ras_n;
output 	[0:0] afi_rst_n;
output 	[0:0] afi_we_n;
output 	[19:0] afi_addr;
output 	[2:0] afi_ba;
output 	[1:0] afi_cke;
output 	[1:0] afi_cs_n;
output 	[9:0] afi_dm;
output 	[4:0] afi_dqs_burst;
output 	[1:0] afi_odt;
output 	[4:0] afi_rdata_en;
output 	[4:0] afi_rdata_en_full;
output 	[79:0] afi_wdata;
output 	[4:0] afi_wdata_valid;
output 	[7:0] cfg_addlat;
output 	[7:0] cfg_bankaddrwidth;
output 	[7:0] cfg_caswrlat;
output 	[7:0] cfg_coladdrwidth;
output 	[7:0] cfg_csaddrwidth;
output 	[7:0] cfg_devicewidth;
output 	[7:0] cfg_interfacewidth;
output 	[7:0] cfg_rowaddrwidth;
output 	[7:0] cfg_tcl;
output 	[7:0] cfg_tmrd;
output 	[15:0] cfg_trefi;
output 	[7:0] cfg_trfc;
output 	[7:0] cfg_twr;
output 	[0:0] afi_mem_clk_disable;
output 	[23:0] cfg_dramconfig;
input 	ctl_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [19:0] hmc_inst_AFIADDR_bus;
wire [2:0] hmc_inst_AFIBA_bus;
wire [1:0] hmc_inst_AFICKE_bus;
wire [1:0] hmc_inst_AFICSN_bus;
wire [9:0] hmc_inst_AFIDM_bus;
wire [4:0] hmc_inst_AFIDQSBURST_bus;
wire [1:0] hmc_inst_AFIODT_bus;
wire [4:0] hmc_inst_AFIRDATAEN_bus;
wire [4:0] hmc_inst_AFIRDATAENFULL_bus;
wire [79:0] hmc_inst_AFIWDATA_bus;
wire [4:0] hmc_inst_AFIWDATAVALID_bus;
wire [4:0] hmc_inst_CFGADDLAT_bus;
wire [2:0] hmc_inst_CFGBANKADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGCASWRLAT_bus;
wire [4:0] hmc_inst_CFGCOLADDRWIDTH_bus;
wire [2:0] hmc_inst_CFGCSADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGDEVICEWIDTH_bus;
wire [7:0] hmc_inst_CFGINTERFACEWIDTH_bus;
wire [4:0] hmc_inst_CFGROWADDRWIDTH_bus;
wire [4:0] hmc_inst_CFGTCL_bus;
wire [3:0] hmc_inst_CFGTMRD_bus;
wire [12:0] hmc_inst_CFGTREFI_bus;
wire [7:0] hmc_inst_CFGTRFC_bus;
wire [3:0] hmc_inst_CFGTWR_bus;
wire [1:0] hmc_inst_CTLMEMCLKDISABLE_bus;
wire [20:0] hmc_inst_DRAMCONFIG_bus;

assign afi_addr[0] = hmc_inst_AFIADDR_bus[0];
assign afi_addr[1] = hmc_inst_AFIADDR_bus[1];
assign afi_addr[2] = hmc_inst_AFIADDR_bus[2];
assign afi_addr[3] = hmc_inst_AFIADDR_bus[3];
assign afi_addr[4] = hmc_inst_AFIADDR_bus[4];
assign afi_addr[5] = hmc_inst_AFIADDR_bus[5];
assign afi_addr[6] = hmc_inst_AFIADDR_bus[6];
assign afi_addr[7] = hmc_inst_AFIADDR_bus[7];
assign afi_addr[8] = hmc_inst_AFIADDR_bus[8];
assign afi_addr[9] = hmc_inst_AFIADDR_bus[9];
assign afi_addr[10] = hmc_inst_AFIADDR_bus[10];
assign afi_addr[11] = hmc_inst_AFIADDR_bus[11];
assign afi_addr[12] = hmc_inst_AFIADDR_bus[12];
assign afi_addr[13] = hmc_inst_AFIADDR_bus[13];
assign afi_addr[14] = hmc_inst_AFIADDR_bus[14];
assign afi_addr[15] = hmc_inst_AFIADDR_bus[15];
assign afi_addr[16] = hmc_inst_AFIADDR_bus[16];
assign afi_addr[17] = hmc_inst_AFIADDR_bus[17];
assign afi_addr[18] = hmc_inst_AFIADDR_bus[18];
assign afi_addr[19] = hmc_inst_AFIADDR_bus[19];

assign afi_ba[0] = hmc_inst_AFIBA_bus[0];
assign afi_ba[1] = hmc_inst_AFIBA_bus[1];
assign afi_ba[2] = hmc_inst_AFIBA_bus[2];

assign afi_cke[0] = hmc_inst_AFICKE_bus[0];
assign afi_cke[1] = hmc_inst_AFICKE_bus[1];

assign afi_cs_n[0] = hmc_inst_AFICSN_bus[0];
assign afi_cs_n[1] = hmc_inst_AFICSN_bus[1];

assign afi_dm[0] = hmc_inst_AFIDM_bus[0];
assign afi_dm[1] = hmc_inst_AFIDM_bus[1];
assign afi_dm[2] = hmc_inst_AFIDM_bus[2];
assign afi_dm[3] = hmc_inst_AFIDM_bus[3];
assign afi_dm[4] = hmc_inst_AFIDM_bus[4];
assign afi_dm[5] = hmc_inst_AFIDM_bus[5];
assign afi_dm[6] = hmc_inst_AFIDM_bus[6];
assign afi_dm[7] = hmc_inst_AFIDM_bus[7];
assign afi_dm[8] = hmc_inst_AFIDM_bus[8];
assign afi_dm[9] = hmc_inst_AFIDM_bus[9];

assign afi_dqs_burst[0] = hmc_inst_AFIDQSBURST_bus[0];
assign afi_dqs_burst[1] = hmc_inst_AFIDQSBURST_bus[1];
assign afi_dqs_burst[2] = hmc_inst_AFIDQSBURST_bus[2];
assign afi_dqs_burst[3] = hmc_inst_AFIDQSBURST_bus[3];
assign afi_dqs_burst[4] = hmc_inst_AFIDQSBURST_bus[4];

assign afi_odt[0] = hmc_inst_AFIODT_bus[0];
assign afi_odt[1] = hmc_inst_AFIODT_bus[1];

assign afi_rdata_en[0] = hmc_inst_AFIRDATAEN_bus[0];
assign afi_rdata_en[1] = hmc_inst_AFIRDATAEN_bus[1];
assign afi_rdata_en[2] = hmc_inst_AFIRDATAEN_bus[2];
assign afi_rdata_en[3] = hmc_inst_AFIRDATAEN_bus[3];
assign afi_rdata_en[4] = hmc_inst_AFIRDATAEN_bus[4];

assign afi_rdata_en_full[0] = hmc_inst_AFIRDATAENFULL_bus[0];
assign afi_rdata_en_full[1] = hmc_inst_AFIRDATAENFULL_bus[1];
assign afi_rdata_en_full[2] = hmc_inst_AFIRDATAENFULL_bus[2];
assign afi_rdata_en_full[3] = hmc_inst_AFIRDATAENFULL_bus[3];
assign afi_rdata_en_full[4] = hmc_inst_AFIRDATAENFULL_bus[4];

assign afi_wdata[0] = hmc_inst_AFIWDATA_bus[0];
assign afi_wdata[1] = hmc_inst_AFIWDATA_bus[1];
assign afi_wdata[2] = hmc_inst_AFIWDATA_bus[2];
assign afi_wdata[3] = hmc_inst_AFIWDATA_bus[3];
assign afi_wdata[4] = hmc_inst_AFIWDATA_bus[4];
assign afi_wdata[5] = hmc_inst_AFIWDATA_bus[5];
assign afi_wdata[6] = hmc_inst_AFIWDATA_bus[6];
assign afi_wdata[7] = hmc_inst_AFIWDATA_bus[7];
assign afi_wdata[8] = hmc_inst_AFIWDATA_bus[8];
assign afi_wdata[9] = hmc_inst_AFIWDATA_bus[9];
assign afi_wdata[10] = hmc_inst_AFIWDATA_bus[10];
assign afi_wdata[11] = hmc_inst_AFIWDATA_bus[11];
assign afi_wdata[12] = hmc_inst_AFIWDATA_bus[12];
assign afi_wdata[13] = hmc_inst_AFIWDATA_bus[13];
assign afi_wdata[14] = hmc_inst_AFIWDATA_bus[14];
assign afi_wdata[15] = hmc_inst_AFIWDATA_bus[15];
assign afi_wdata[16] = hmc_inst_AFIWDATA_bus[16];
assign afi_wdata[17] = hmc_inst_AFIWDATA_bus[17];
assign afi_wdata[18] = hmc_inst_AFIWDATA_bus[18];
assign afi_wdata[19] = hmc_inst_AFIWDATA_bus[19];
assign afi_wdata[20] = hmc_inst_AFIWDATA_bus[20];
assign afi_wdata[21] = hmc_inst_AFIWDATA_bus[21];
assign afi_wdata[22] = hmc_inst_AFIWDATA_bus[22];
assign afi_wdata[23] = hmc_inst_AFIWDATA_bus[23];
assign afi_wdata[24] = hmc_inst_AFIWDATA_bus[24];
assign afi_wdata[25] = hmc_inst_AFIWDATA_bus[25];
assign afi_wdata[26] = hmc_inst_AFIWDATA_bus[26];
assign afi_wdata[27] = hmc_inst_AFIWDATA_bus[27];
assign afi_wdata[28] = hmc_inst_AFIWDATA_bus[28];
assign afi_wdata[29] = hmc_inst_AFIWDATA_bus[29];
assign afi_wdata[30] = hmc_inst_AFIWDATA_bus[30];
assign afi_wdata[31] = hmc_inst_AFIWDATA_bus[31];
assign afi_wdata[32] = hmc_inst_AFIWDATA_bus[32];
assign afi_wdata[33] = hmc_inst_AFIWDATA_bus[33];
assign afi_wdata[34] = hmc_inst_AFIWDATA_bus[34];
assign afi_wdata[35] = hmc_inst_AFIWDATA_bus[35];
assign afi_wdata[36] = hmc_inst_AFIWDATA_bus[36];
assign afi_wdata[37] = hmc_inst_AFIWDATA_bus[37];
assign afi_wdata[38] = hmc_inst_AFIWDATA_bus[38];
assign afi_wdata[39] = hmc_inst_AFIWDATA_bus[39];
assign afi_wdata[40] = hmc_inst_AFIWDATA_bus[40];
assign afi_wdata[41] = hmc_inst_AFIWDATA_bus[41];
assign afi_wdata[42] = hmc_inst_AFIWDATA_bus[42];
assign afi_wdata[43] = hmc_inst_AFIWDATA_bus[43];
assign afi_wdata[44] = hmc_inst_AFIWDATA_bus[44];
assign afi_wdata[45] = hmc_inst_AFIWDATA_bus[45];
assign afi_wdata[46] = hmc_inst_AFIWDATA_bus[46];
assign afi_wdata[47] = hmc_inst_AFIWDATA_bus[47];
assign afi_wdata[48] = hmc_inst_AFIWDATA_bus[48];
assign afi_wdata[49] = hmc_inst_AFIWDATA_bus[49];
assign afi_wdata[50] = hmc_inst_AFIWDATA_bus[50];
assign afi_wdata[51] = hmc_inst_AFIWDATA_bus[51];
assign afi_wdata[52] = hmc_inst_AFIWDATA_bus[52];
assign afi_wdata[53] = hmc_inst_AFIWDATA_bus[53];
assign afi_wdata[54] = hmc_inst_AFIWDATA_bus[54];
assign afi_wdata[55] = hmc_inst_AFIWDATA_bus[55];
assign afi_wdata[56] = hmc_inst_AFIWDATA_bus[56];
assign afi_wdata[57] = hmc_inst_AFIWDATA_bus[57];
assign afi_wdata[58] = hmc_inst_AFIWDATA_bus[58];
assign afi_wdata[59] = hmc_inst_AFIWDATA_bus[59];
assign afi_wdata[60] = hmc_inst_AFIWDATA_bus[60];
assign afi_wdata[61] = hmc_inst_AFIWDATA_bus[61];
assign afi_wdata[62] = hmc_inst_AFIWDATA_bus[62];
assign afi_wdata[63] = hmc_inst_AFIWDATA_bus[63];
assign afi_wdata[64] = hmc_inst_AFIWDATA_bus[64];
assign afi_wdata[65] = hmc_inst_AFIWDATA_bus[65];
assign afi_wdata[66] = hmc_inst_AFIWDATA_bus[66];
assign afi_wdata[67] = hmc_inst_AFIWDATA_bus[67];
assign afi_wdata[68] = hmc_inst_AFIWDATA_bus[68];
assign afi_wdata[69] = hmc_inst_AFIWDATA_bus[69];
assign afi_wdata[70] = hmc_inst_AFIWDATA_bus[70];
assign afi_wdata[71] = hmc_inst_AFIWDATA_bus[71];
assign afi_wdata[72] = hmc_inst_AFIWDATA_bus[72];
assign afi_wdata[73] = hmc_inst_AFIWDATA_bus[73];
assign afi_wdata[74] = hmc_inst_AFIWDATA_bus[74];
assign afi_wdata[75] = hmc_inst_AFIWDATA_bus[75];
assign afi_wdata[76] = hmc_inst_AFIWDATA_bus[76];
assign afi_wdata[77] = hmc_inst_AFIWDATA_bus[77];
assign afi_wdata[78] = hmc_inst_AFIWDATA_bus[78];
assign afi_wdata[79] = hmc_inst_AFIWDATA_bus[79];

assign afi_wdata_valid[0] = hmc_inst_AFIWDATAVALID_bus[0];
assign afi_wdata_valid[1] = hmc_inst_AFIWDATAVALID_bus[1];
assign afi_wdata_valid[2] = hmc_inst_AFIWDATAVALID_bus[2];
assign afi_wdata_valid[3] = hmc_inst_AFIWDATAVALID_bus[3];
assign afi_wdata_valid[4] = hmc_inst_AFIWDATAVALID_bus[4];

assign cfg_addlat[0] = hmc_inst_CFGADDLAT_bus[0];
assign cfg_addlat[1] = hmc_inst_CFGADDLAT_bus[1];
assign cfg_addlat[2] = hmc_inst_CFGADDLAT_bus[2];
assign cfg_addlat[3] = hmc_inst_CFGADDLAT_bus[3];
assign cfg_addlat[4] = hmc_inst_CFGADDLAT_bus[4];

assign cfg_bankaddrwidth[0] = hmc_inst_CFGBANKADDRWIDTH_bus[0];
assign cfg_bankaddrwidth[1] = hmc_inst_CFGBANKADDRWIDTH_bus[1];
assign cfg_bankaddrwidth[2] = hmc_inst_CFGBANKADDRWIDTH_bus[2];

assign cfg_caswrlat[0] = hmc_inst_CFGCASWRLAT_bus[0];
assign cfg_caswrlat[1] = hmc_inst_CFGCASWRLAT_bus[1];
assign cfg_caswrlat[2] = hmc_inst_CFGCASWRLAT_bus[2];
assign cfg_caswrlat[3] = hmc_inst_CFGCASWRLAT_bus[3];

assign cfg_coladdrwidth[0] = hmc_inst_CFGCOLADDRWIDTH_bus[0];
assign cfg_coladdrwidth[1] = hmc_inst_CFGCOLADDRWIDTH_bus[1];
assign cfg_coladdrwidth[2] = hmc_inst_CFGCOLADDRWIDTH_bus[2];
assign cfg_coladdrwidth[3] = hmc_inst_CFGCOLADDRWIDTH_bus[3];
assign cfg_coladdrwidth[4] = hmc_inst_CFGCOLADDRWIDTH_bus[4];

assign cfg_csaddrwidth[0] = hmc_inst_CFGCSADDRWIDTH_bus[0];
assign cfg_csaddrwidth[1] = hmc_inst_CFGCSADDRWIDTH_bus[1];
assign cfg_csaddrwidth[2] = hmc_inst_CFGCSADDRWIDTH_bus[2];

assign cfg_devicewidth[0] = hmc_inst_CFGDEVICEWIDTH_bus[0];
assign cfg_devicewidth[1] = hmc_inst_CFGDEVICEWIDTH_bus[1];
assign cfg_devicewidth[2] = hmc_inst_CFGDEVICEWIDTH_bus[2];
assign cfg_devicewidth[3] = hmc_inst_CFGDEVICEWIDTH_bus[3];

assign cfg_interfacewidth[0] = hmc_inst_CFGINTERFACEWIDTH_bus[0];
assign cfg_interfacewidth[1] = hmc_inst_CFGINTERFACEWIDTH_bus[1];
assign cfg_interfacewidth[2] = hmc_inst_CFGINTERFACEWIDTH_bus[2];
assign cfg_interfacewidth[3] = hmc_inst_CFGINTERFACEWIDTH_bus[3];
assign cfg_interfacewidth[4] = hmc_inst_CFGINTERFACEWIDTH_bus[4];
assign cfg_interfacewidth[5] = hmc_inst_CFGINTERFACEWIDTH_bus[5];
assign cfg_interfacewidth[6] = hmc_inst_CFGINTERFACEWIDTH_bus[6];
assign cfg_interfacewidth[7] = hmc_inst_CFGINTERFACEWIDTH_bus[7];

assign cfg_rowaddrwidth[0] = hmc_inst_CFGROWADDRWIDTH_bus[0];
assign cfg_rowaddrwidth[1] = hmc_inst_CFGROWADDRWIDTH_bus[1];
assign cfg_rowaddrwidth[2] = hmc_inst_CFGROWADDRWIDTH_bus[2];
assign cfg_rowaddrwidth[3] = hmc_inst_CFGROWADDRWIDTH_bus[3];
assign cfg_rowaddrwidth[4] = hmc_inst_CFGROWADDRWIDTH_bus[4];

assign cfg_tcl[0] = hmc_inst_CFGTCL_bus[0];
assign cfg_tcl[1] = hmc_inst_CFGTCL_bus[1];
assign cfg_tcl[2] = hmc_inst_CFGTCL_bus[2];
assign cfg_tcl[3] = hmc_inst_CFGTCL_bus[3];
assign cfg_tcl[4] = hmc_inst_CFGTCL_bus[4];

assign cfg_tmrd[0] = hmc_inst_CFGTMRD_bus[0];
assign cfg_tmrd[1] = hmc_inst_CFGTMRD_bus[1];
assign cfg_tmrd[2] = hmc_inst_CFGTMRD_bus[2];
assign cfg_tmrd[3] = hmc_inst_CFGTMRD_bus[3];

assign cfg_trefi[0] = hmc_inst_CFGTREFI_bus[0];
assign cfg_trefi[1] = hmc_inst_CFGTREFI_bus[1];
assign cfg_trefi[2] = hmc_inst_CFGTREFI_bus[2];
assign cfg_trefi[3] = hmc_inst_CFGTREFI_bus[3];
assign cfg_trefi[4] = hmc_inst_CFGTREFI_bus[4];
assign cfg_trefi[5] = hmc_inst_CFGTREFI_bus[5];
assign cfg_trefi[6] = hmc_inst_CFGTREFI_bus[6];
assign cfg_trefi[7] = hmc_inst_CFGTREFI_bus[7];
assign cfg_trefi[8] = hmc_inst_CFGTREFI_bus[8];
assign cfg_trefi[9] = hmc_inst_CFGTREFI_bus[9];
assign cfg_trefi[10] = hmc_inst_CFGTREFI_bus[10];
assign cfg_trefi[11] = hmc_inst_CFGTREFI_bus[11];
assign cfg_trefi[12] = hmc_inst_CFGTREFI_bus[12];

assign cfg_trfc[0] = hmc_inst_CFGTRFC_bus[0];
assign cfg_trfc[1] = hmc_inst_CFGTRFC_bus[1];
assign cfg_trfc[2] = hmc_inst_CFGTRFC_bus[2];
assign cfg_trfc[3] = hmc_inst_CFGTRFC_bus[3];
assign cfg_trfc[4] = hmc_inst_CFGTRFC_bus[4];
assign cfg_trfc[5] = hmc_inst_CFGTRFC_bus[5];
assign cfg_trfc[6] = hmc_inst_CFGTRFC_bus[6];
assign cfg_trfc[7] = hmc_inst_CFGTRFC_bus[7];

assign cfg_twr[0] = hmc_inst_CFGTWR_bus[0];
assign cfg_twr[1] = hmc_inst_CFGTWR_bus[1];
assign cfg_twr[2] = hmc_inst_CFGTWR_bus[2];
assign cfg_twr[3] = hmc_inst_CFGTWR_bus[3];

assign afi_mem_clk_disable[0] = hmc_inst_CTLMEMCLKDISABLE_bus[0];

assign cfg_dramconfig[0] = hmc_inst_DRAMCONFIG_bus[0];
assign cfg_dramconfig[1] = hmc_inst_DRAMCONFIG_bus[1];
assign cfg_dramconfig[2] = hmc_inst_DRAMCONFIG_bus[2];
assign cfg_dramconfig[3] = hmc_inst_DRAMCONFIG_bus[3];
assign cfg_dramconfig[4] = hmc_inst_DRAMCONFIG_bus[4];
assign cfg_dramconfig[5] = hmc_inst_DRAMCONFIG_bus[5];
assign cfg_dramconfig[6] = hmc_inst_DRAMCONFIG_bus[6];
assign cfg_dramconfig[7] = hmc_inst_DRAMCONFIG_bus[7];
assign cfg_dramconfig[8] = hmc_inst_DRAMCONFIG_bus[8];
assign cfg_dramconfig[9] = hmc_inst_DRAMCONFIG_bus[9];
assign cfg_dramconfig[10] = hmc_inst_DRAMCONFIG_bus[10];
assign cfg_dramconfig[11] = hmc_inst_DRAMCONFIG_bus[11];
assign cfg_dramconfig[12] = hmc_inst_DRAMCONFIG_bus[12];
assign cfg_dramconfig[13] = hmc_inst_DRAMCONFIG_bus[13];
assign cfg_dramconfig[14] = hmc_inst_DRAMCONFIG_bus[14];
assign cfg_dramconfig[15] = hmc_inst_DRAMCONFIG_bus[15];
assign cfg_dramconfig[16] = hmc_inst_DRAMCONFIG_bus[16];
assign cfg_dramconfig[17] = hmc_inst_DRAMCONFIG_bus[17];
assign cfg_dramconfig[18] = hmc_inst_DRAMCONFIG_bus[18];
assign cfg_dramconfig[19] = hmc_inst_DRAMCONFIG_bus[19];
assign cfg_dramconfig[20] = hmc_inst_DRAMCONFIG_bus[20];

cyclonev_hmc hmc_inst(
	.afirdatavalid(afi_rdata_valid[0]),
	.csrclk(gnd),
	.csrdin(gnd),
	.csren(gnd),
	.ctlcalfail(afi_cal_fail),
	.ctlcalsuccess(afi_cal_success),
	.ctlclk(ctl_clk),
	.ctlresetn(ctl_reset_n),
	.globalresetn(gnd),
	.iavstcmdresetn0(vcc),
	.iavstcmdresetn1(vcc),
	.iavstcmdresetn2(vcc),
	.iavstcmdresetn3(vcc),
	.iavstcmdresetn4(vcc),
	.iavstcmdresetn5(vcc),
	.iavstrdclk0(gnd),
	.iavstrdclk1(gnd),
	.iavstrdclk2(gnd),
	.iavstrdclk3(gnd),
	.iavstrdready0(vcc),
	.iavstrdready1(vcc),
	.iavstrdready2(vcc),
	.iavstrdready3(vcc),
	.iavstrdresetn0(vcc),
	.iavstrdresetn1(vcc),
	.iavstrdresetn2(vcc),
	.iavstrdresetn3(vcc),
	.iavstwrackready0(vcc),
	.iavstwrackready1(vcc),
	.iavstwrackready2(vcc),
	.iavstwrackready3(vcc),
	.iavstwrackready4(vcc),
	.iavstwrackready5(vcc),
	.iavstwrclk0(gnd),
	.iavstwrclk1(gnd),
	.iavstwrclk2(gnd),
	.iavstwrclk3(gnd),
	.iavstwrresetn0(vcc),
	.iavstwrresetn1(vcc),
	.iavstwrresetn2(vcc),
	.iavstwrresetn3(vcc),
	.localdeeppowerdnreq(gnd),
	.localrefreshreq(gnd),
	.localselfrfshreq(gnd),
	.mmrbe(gnd),
	.mmrburstbegin(vcc),
	.mmrclk(gnd),
	.mmrreadreq(gnd),
	.mmrresetn(vcc),
	.mmrwritereq(gnd),
	.portclk0(gnd),
	.portclk1(gnd),
	.portclk2(gnd),
	.portclk3(gnd),
	.portclk4(gnd),
	.portclk5(gnd),
	.scanenable(gnd),
	.scbe(gnd),
	.scburstbegin(gnd),
	.scclk(gnd),
	.screadreq(gnd),
	.scresetn(vcc),
	.scwritereq(gnd),
	.afirdata({afi_rdata[79],afi_rdata[78],afi_rdata[77],afi_rdata[76],afi_rdata[75],afi_rdata[74],afi_rdata[73],afi_rdata[72],afi_rdata[71],afi_rdata[70],afi_rdata[69],afi_rdata[68],afi_rdata[67],afi_rdata[66],afi_rdata[65],afi_rdata[64],afi_rdata[63],afi_rdata[62],afi_rdata[61],afi_rdata[60],afi_rdata[59],afi_rdata[58],afi_rdata[57],afi_rdata[56],afi_rdata[55],afi_rdata[54],afi_rdata[53],afi_rdata[52],
afi_rdata[51],afi_rdata[50],afi_rdata[49],afi_rdata[48],afi_rdata[47],afi_rdata[46],afi_rdata[45],afi_rdata[44],afi_rdata[43],afi_rdata[42],afi_rdata[41],afi_rdata[40],afi_rdata[39],afi_rdata[38],afi_rdata[37],afi_rdata[36],afi_rdata[35],afi_rdata[34],afi_rdata[33],afi_rdata[32],afi_rdata[31],afi_rdata[30],afi_rdata[29],afi_rdata[28],afi_rdata[27],afi_rdata[26],afi_rdata[25],afi_rdata[24],
afi_rdata[23],afi_rdata[22],afi_rdata[21],afi_rdata[20],afi_rdata[19],afi_rdata[18],afi_rdata[17],afi_rdata[16],afi_rdata[15],afi_rdata[14],afi_rdata[13],afi_rdata[12],afi_rdata[11],afi_rdata[10],afi_rdata[9],afi_rdata[8],afi_rdata[7],afi_rdata[6],afi_rdata[5],afi_rdata[4],afi_rdata[3],afi_rdata[2],afi_rdata[1],afi_rdata[0]}),
	.afiseqbusy({gnd,gnd}),
	.afiwlat({afi_wlat[3],afi_wlat[2],afi_wlat[1],afi_wlat[0]}),
	.bondingin1({gnd,gnd,gnd,gnd}),
	.bondingin2({gnd,gnd,gnd,gnd,gnd,gnd}),
	.bondingin3({gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata4({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata5({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.localdeeppowerdnchip({gnd,gnd}),
	.localrefreshchip({gnd,gnd}),
	.localselfrfshchip({gnd,gnd}),
	.mmraddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.mmrburstcount({gnd,vcc}),
	.mmrwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scburstcount({gnd,gnd}),
	.scwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.aficasn(afi_cas_n[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.csrdout(),
	.ctlcalreq(),
	.ctlinitreq(),
	.localdeeppowerdnack(),
	.localinitdone(),
	.localpowerdownack(),
	.localrefreshack(),
	.localselfrfshack(),
	.localstsctlempty(),
	.mmrrdatavalid(),
	.mmrwaitrequest(),
	.oammready0(),
	.oammready1(),
	.oammready2(),
	.oammready3(),
	.oammready4(),
	.oammready5(),
	.ordavstvalid0(),
	.ordavstvalid1(),
	.ordavstvalid2(),
	.ordavstvalid3(),
	.owrackavstdata0(),
	.owrackavstdata1(),
	.owrackavstdata2(),
	.owrackavstdata3(),
	.owrackavstdata4(),
	.owrackavstdata5(),
	.owrackavstvalid0(),
	.owrackavstvalid1(),
	.owrackavstvalid2(),
	.owrackavstvalid3(),
	.owrackavstvalid4(),
	.owrackavstvalid5(),
	.scrdatavalid(),
	.scwaitrequest(),
	.afiaddr(hmc_inst_AFIADDR_bus),
	.afiba(hmc_inst_AFIBA_bus),
	.aficke(hmc_inst_AFICKE_bus),
	.aficsn(hmc_inst_AFICSN_bus),
	.afictllongidle(),
	.afictlrefreshdone(),
	.afidm(hmc_inst_AFIDM_bus),
	.afidqsburst(hmc_inst_AFIDQSBURST_bus),
	.afiodt(hmc_inst_AFIODT_bus),
	.afirdataen(hmc_inst_AFIRDATAEN_bus),
	.afirdataenfull(hmc_inst_AFIRDATAENFULL_bus),
	.afiwdata(hmc_inst_AFIWDATA_bus),
	.afiwdatavalid(hmc_inst_AFIWDATAVALID_bus),
	.bondingout1(),
	.bondingout2(),
	.bondingout3(),
	.cfgaddlat(hmc_inst_CFGADDLAT_bus),
	.cfgbankaddrwidth(hmc_inst_CFGBANKADDRWIDTH_bus),
	.cfgcaswrlat(hmc_inst_CFGCASWRLAT_bus),
	.cfgcoladdrwidth(hmc_inst_CFGCOLADDRWIDTH_bus),
	.cfgcsaddrwidth(hmc_inst_CFGCSADDRWIDTH_bus),
	.cfgdevicewidth(hmc_inst_CFGDEVICEWIDTH_bus),
	.cfginterfacewidth(hmc_inst_CFGINTERFACEWIDTH_bus),
	.cfgrowaddrwidth(hmc_inst_CFGROWADDRWIDTH_bus),
	.cfgtcl(hmc_inst_CFGTCL_bus),
	.cfgtmrd(hmc_inst_CFGTMRD_bus),
	.cfgtrefi(hmc_inst_CFGTREFI_bus),
	.cfgtrfc(hmc_inst_CFGTRFC_bus),
	.cfgtwr(hmc_inst_CFGTWR_bus),
	.ctlcalbytelaneseln(),
	.ctlmemclkdisable(hmc_inst_CTLMEMCLKDISABLE_bus),
	.dramconfig(hmc_inst_DRAMCONFIG_bus),
	.mmrrdata(),
	.ordavstdata0(),
	.ordavstdata1(),
	.ordavstdata2(),
	.ordavstdata3(),
	.scrdata());
defparam hmc_inst.attr_counter_one_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_reset = "disabled";
defparam hmc_inst.attr_counter_zero_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_reset = "disabled";
defparam hmc_inst.attr_debug_select_byte = 32'b00000000000000000000000000000000;
defparam hmc_inst.attr_static_config_valid = "disabled";
defparam hmc_inst.auto_pch_enable_0 = "disabled";
defparam hmc_inst.auto_pch_enable_1 = "disabled";
defparam hmc_inst.auto_pch_enable_2 = "disabled";
defparam hmc_inst.auto_pch_enable_3 = "disabled";
defparam hmc_inst.auto_pch_enable_4 = "disabled";
defparam hmc_inst.auto_pch_enable_5 = "disabled";
defparam hmc_inst.cal_req = "disabled";
defparam hmc_inst.cfg_burst_length = "bl_8";
defparam hmc_inst.cfg_interface_width = "dwidth_32";
defparam hmc_inst.cfg_self_rfsh_exit_cycles = "self_rfsh_exit_cycles_512";
defparam hmc_inst.cfg_starve_limit = "starve_limit_10";
defparam hmc_inst.cfg_type = "ddr3";
defparam hmc_inst.clr_intr = "no_clr_intr";
defparam hmc_inst.cmd_port_in_use_0 = "false";
defparam hmc_inst.cmd_port_in_use_1 = "false";
defparam hmc_inst.cmd_port_in_use_2 = "false";
defparam hmc_inst.cmd_port_in_use_3 = "false";
defparam hmc_inst.cmd_port_in_use_4 = "false";
defparam hmc_inst.cmd_port_in_use_5 = "false";
defparam hmc_inst.cport0_rdy_almost_full = "not_full";
defparam hmc_inst.cport0_rfifo_map = "fifo_0";
defparam hmc_inst.cport0_type = "disable";
defparam hmc_inst.cport0_wfifo_map = "fifo_0";
defparam hmc_inst.cport1_rdy_almost_full = "not_full";
defparam hmc_inst.cport1_rfifo_map = "fifo_0";
defparam hmc_inst.cport1_type = "disable";
defparam hmc_inst.cport1_wfifo_map = "fifo_0";
defparam hmc_inst.cport2_rdy_almost_full = "not_full";
defparam hmc_inst.cport2_rfifo_map = "fifo_0";
defparam hmc_inst.cport2_type = "disable";
defparam hmc_inst.cport2_wfifo_map = "fifo_0";
defparam hmc_inst.cport3_rdy_almost_full = "not_full";
defparam hmc_inst.cport3_rfifo_map = "fifo_0";
defparam hmc_inst.cport3_type = "disable";
defparam hmc_inst.cport3_wfifo_map = "fifo_0";
defparam hmc_inst.cport4_rdy_almost_full = "not_full";
defparam hmc_inst.cport4_rfifo_map = "fifo_0";
defparam hmc_inst.cport4_type = "disable";
defparam hmc_inst.cport4_wfifo_map = "fifo_0";
defparam hmc_inst.cport5_rdy_almost_full = "not_full";
defparam hmc_inst.cport5_rfifo_map = "fifo_0";
defparam hmc_inst.cport5_type = "disable";
defparam hmc_inst.cport5_wfifo_map = "fifo_0";
defparam hmc_inst.ctl_addr_order = "chip_row_bank_col";
defparam hmc_inst.ctl_ecc_enabled = "ctl_ecc_disabled";
defparam hmc_inst.ctl_ecc_rmw_enabled = "ctl_ecc_rmw_disabled";
defparam hmc_inst.ctl_regdimm_enabled = "regdimm_disabled";
defparam hmc_inst.ctl_usr_refresh = "ctl_usr_refresh_disabled";
defparam hmc_inst.ctrl_width = "data_width_64_bit";
defparam hmc_inst.cyc_to_rld_jars_0 = 1;
defparam hmc_inst.cyc_to_rld_jars_1 = 1;
defparam hmc_inst.cyc_to_rld_jars_2 = 1;
defparam hmc_inst.cyc_to_rld_jars_3 = 1;
defparam hmc_inst.cyc_to_rld_jars_4 = 1;
defparam hmc_inst.cyc_to_rld_jars_5 = 1;
defparam hmc_inst.delay_bonding = "bonding_latency_0";
defparam hmc_inst.dfx_bypass_enable = "dfx_bypass_disabled";
defparam hmc_inst.disable_merging = "merging_enabled";
defparam hmc_inst.ecc_dq_width = "ecc_dq_width_0";
defparam hmc_inst.enable_atpg = "disabled";
defparam hmc_inst.enable_bonding_0 = "disabled";
defparam hmc_inst.enable_bonding_1 = "disabled";
defparam hmc_inst.enable_bonding_2 = "disabled";
defparam hmc_inst.enable_bonding_3 = "disabled";
defparam hmc_inst.enable_bonding_4 = "disabled";
defparam hmc_inst.enable_bonding_5 = "disabled";
defparam hmc_inst.enable_bonding_wrapback = "disabled";
defparam hmc_inst.enable_burst_interrupt = "disabled";
defparam hmc_inst.enable_burst_terminate = "disabled";
defparam hmc_inst.enable_dqs_tracking = "enabled";
defparam hmc_inst.enable_ecc_code_overwrites = "disabled";
defparam hmc_inst.enable_fast_exit_ppd = "disabled";
defparam hmc_inst.enable_intr = "disabled";
defparam hmc_inst.enable_no_dm = "disabled";
defparam hmc_inst.enable_pipelineglobal = "disabled";
defparam hmc_inst.extra_ctl_clk_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_act_to_act_diff_bank = 0;
defparam hmc_inst.extra_ctl_clk_act_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_act_to_rdwr = 0;
defparam hmc_inst.extra_ctl_clk_arf_period = 0;
defparam hmc_inst.extra_ctl_clk_arf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_four_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_pch_all_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pch_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pdn_period = 0;
defparam hmc_inst.extra_ctl_clk_pdn_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd_diff_chip = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_wr = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_bc = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_diff_chip = 2;
defparam hmc_inst.extra_ctl_clk_srf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_srf_to_zq_cal = 0;
defparam hmc_inst.extra_ctl_clk_wr_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_rd = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_bc = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_diff_chip = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_wr = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_wr_diff_chip = 0;
defparam hmc_inst.gen_dbe = "gen_dbe_disabled";
defparam hmc_inst.gen_sbe = "gen_sbe_disabled";
defparam hmc_inst.inc_sync = "fifo_set_2";
defparam hmc_inst.local_if_cs_width = "addr_width_0";
defparam hmc_inst.mask_corr_dropped_intr = "disabled";
defparam hmc_inst.mask_dbe_intr = "disabled";
defparam hmc_inst.mask_sbe_intr = "disabled";
defparam hmc_inst.mem_auto_pd_cycles = 0;
defparam hmc_inst.mem_clk_entry_cycles = 10;
defparam hmc_inst.mem_if_al = "al_0";
defparam hmc_inst.mem_if_bankaddr_width = "addr_width_3";
defparam hmc_inst.mem_if_burstlength = "mem_if_burstlength_8";
defparam hmc_inst.mem_if_coladdr_width = "addr_width_10";
defparam hmc_inst.mem_if_cs_per_rank = "mem_if_cs_per_rank_1";
defparam hmc_inst.mem_if_cs_width = "mem_if_cs_width_1";
defparam hmc_inst.mem_if_dq_per_chip = "mem_if_dq_per_chip_8";
defparam hmc_inst.mem_if_dqs_width = "dqs_width_4";
defparam hmc_inst.mem_if_dwidth = "mem_if_dwidth_32";
defparam hmc_inst.mem_if_memtype = "ddr3_sdram";
defparam hmc_inst.mem_if_rowaddr_width = "addr_width_15";
defparam hmc_inst.mem_if_speedbin = "ddr3_1600_8_8_8";
defparam hmc_inst.mem_if_tccd = "tccd_4";
defparam hmc_inst.mem_if_tcl = "tcl_11";
defparam hmc_inst.mem_if_tcwl = "tcwl_8";
defparam hmc_inst.mem_if_tfaw = "tfaw_12";
defparam hmc_inst.mem_if_tmrd = "tmrd_4";
defparam hmc_inst.mem_if_tras = "tras_14";
defparam hmc_inst.mem_if_trc = "trc_20";
defparam hmc_inst.mem_if_trcd = "trcd_6";
defparam hmc_inst.mem_if_trefi = 3120;
defparam hmc_inst.mem_if_trfc = 104;
defparam hmc_inst.mem_if_trp = "trp_6";
defparam hmc_inst.mem_if_trrd = "trrd_3";
defparam hmc_inst.mem_if_trtp = "trtp_3";
defparam hmc_inst.mem_if_twr = "twr_6";
defparam hmc_inst.mem_if_twtr = "twtr_4";
defparam hmc_inst.mmr_cfg_mem_bl = "mp_bl_8";
defparam hmc_inst.output_regd = "disabled";
defparam hmc_inst.pdn_exit_cycles = "slow_exit";
defparam hmc_inst.port0_width = "port_32_bit";
defparam hmc_inst.port1_width = "port_32_bit";
defparam hmc_inst.port2_width = "port_32_bit";
defparam hmc_inst.port3_width = "port_32_bit";
defparam hmc_inst.port4_width = "port_32_bit";
defparam hmc_inst.port5_width = "port_32_bit";
defparam hmc_inst.power_saving_exit_cycles = 5;
defparam hmc_inst.priority_0_0 = "weight_0";
defparam hmc_inst.priority_0_1 = "weight_0";
defparam hmc_inst.priority_0_2 = "weight_0";
defparam hmc_inst.priority_0_3 = "weight_0";
defparam hmc_inst.priority_0_4 = "weight_0";
defparam hmc_inst.priority_0_5 = "weight_0";
defparam hmc_inst.priority_1_0 = "weight_0";
defparam hmc_inst.priority_1_1 = "weight_0";
defparam hmc_inst.priority_1_2 = "weight_0";
defparam hmc_inst.priority_1_3 = "weight_0";
defparam hmc_inst.priority_1_4 = "weight_0";
defparam hmc_inst.priority_1_5 = "weight_0";
defparam hmc_inst.priority_2_0 = "weight_0";
defparam hmc_inst.priority_2_1 = "weight_0";
defparam hmc_inst.priority_2_2 = "weight_0";
defparam hmc_inst.priority_2_3 = "weight_0";
defparam hmc_inst.priority_2_4 = "weight_0";
defparam hmc_inst.priority_2_5 = "weight_0";
defparam hmc_inst.priority_3_0 = "weight_0";
defparam hmc_inst.priority_3_1 = "weight_0";
defparam hmc_inst.priority_3_2 = "weight_0";
defparam hmc_inst.priority_3_3 = "weight_0";
defparam hmc_inst.priority_3_4 = "weight_0";
defparam hmc_inst.priority_3_5 = "weight_0";
defparam hmc_inst.priority_4_0 = "weight_0";
defparam hmc_inst.priority_4_1 = "weight_0";
defparam hmc_inst.priority_4_2 = "weight_0";
defparam hmc_inst.priority_4_3 = "weight_0";
defparam hmc_inst.priority_4_4 = "weight_0";
defparam hmc_inst.priority_4_5 = "weight_0";
defparam hmc_inst.priority_5_0 = "weight_0";
defparam hmc_inst.priority_5_1 = "weight_0";
defparam hmc_inst.priority_5_2 = "weight_0";
defparam hmc_inst.priority_5_3 = "weight_0";
defparam hmc_inst.priority_5_4 = "weight_0";
defparam hmc_inst.priority_5_5 = "weight_0";
defparam hmc_inst.priority_6_0 = "weight_0";
defparam hmc_inst.priority_6_1 = "weight_0";
defparam hmc_inst.priority_6_2 = "weight_0";
defparam hmc_inst.priority_6_3 = "weight_0";
defparam hmc_inst.priority_6_4 = "weight_0";
defparam hmc_inst.priority_6_5 = "weight_0";
defparam hmc_inst.priority_7_0 = "weight_0";
defparam hmc_inst.priority_7_1 = "weight_0";
defparam hmc_inst.priority_7_2 = "weight_0";
defparam hmc_inst.priority_7_3 = "weight_0";
defparam hmc_inst.priority_7_4 = "weight_0";
defparam hmc_inst.priority_7_5 = "weight_0";
defparam hmc_inst.priority_remap = 0;
defparam hmc_inst.rcfg_static_weight_0 = "weight_0";
defparam hmc_inst.rcfg_static_weight_1 = "weight_0";
defparam hmc_inst.rcfg_static_weight_2 = "weight_0";
defparam hmc_inst.rcfg_static_weight_3 = "weight_0";
defparam hmc_inst.rcfg_static_weight_4 = "weight_0";
defparam hmc_inst.rcfg_static_weight_5 = "weight_0";
defparam hmc_inst.rcfg_sum_wt_priority_0 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_1 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_2 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_3 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_4 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_5 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_6 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_7 = 0;
defparam hmc_inst.rcfg_user_priority_0 = "priority_1";
defparam hmc_inst.rcfg_user_priority_1 = "priority_1";
defparam hmc_inst.rcfg_user_priority_2 = "priority_1";
defparam hmc_inst.rcfg_user_priority_3 = "priority_1";
defparam hmc_inst.rcfg_user_priority_4 = "priority_1";
defparam hmc_inst.rcfg_user_priority_5 = "priority_1";
defparam hmc_inst.rd_dwidth_0 = "dwidth_0";
defparam hmc_inst.rd_dwidth_1 = "dwidth_0";
defparam hmc_inst.rd_dwidth_2 = "dwidth_0";
defparam hmc_inst.rd_dwidth_3 = "dwidth_0";
defparam hmc_inst.rd_dwidth_4 = "dwidth_0";
defparam hmc_inst.rd_dwidth_5 = "dwidth_0";
defparam hmc_inst.rd_fifo_in_use_0 = "false";
defparam hmc_inst.rd_fifo_in_use_1 = "false";
defparam hmc_inst.rd_fifo_in_use_2 = "false";
defparam hmc_inst.rd_fifo_in_use_3 = "false";
defparam hmc_inst.rd_port_info_0 = "use_no";
defparam hmc_inst.rd_port_info_1 = "use_no";
defparam hmc_inst.rd_port_info_2 = "use_no";
defparam hmc_inst.rd_port_info_3 = "use_no";
defparam hmc_inst.rd_port_info_4 = "use_no";
defparam hmc_inst.rd_port_info_5 = "use_no";
defparam hmc_inst.read_odt_chip = "odt_disabled";
defparam hmc_inst.reorder_data = "data_reordering";
defparam hmc_inst.rfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.single_ready_0 = "concatenate_rdy";
defparam hmc_inst.single_ready_1 = "concatenate_rdy";
defparam hmc_inst.single_ready_2 = "concatenate_rdy";
defparam hmc_inst.single_ready_3 = "concatenate_rdy";
defparam hmc_inst.static_weight_0 = "weight_0";
defparam hmc_inst.static_weight_1 = "weight_0";
defparam hmc_inst.static_weight_2 = "weight_0";
defparam hmc_inst.static_weight_3 = "weight_0";
defparam hmc_inst.static_weight_4 = "weight_0";
defparam hmc_inst.static_weight_5 = "weight_0";
defparam hmc_inst.sum_wt_priority_0 = 0;
defparam hmc_inst.sum_wt_priority_1 = 0;
defparam hmc_inst.sum_wt_priority_2 = 0;
defparam hmc_inst.sum_wt_priority_3 = 0;
defparam hmc_inst.sum_wt_priority_4 = 0;
defparam hmc_inst.sum_wt_priority_5 = 0;
defparam hmc_inst.sum_wt_priority_6 = 0;
defparam hmc_inst.sum_wt_priority_7 = 0;
defparam hmc_inst.sync_mode_0 = "asynchronous";
defparam hmc_inst.sync_mode_1 = "asynchronous";
defparam hmc_inst.sync_mode_2 = "asynchronous";
defparam hmc_inst.sync_mode_3 = "asynchronous";
defparam hmc_inst.sync_mode_4 = "asynchronous";
defparam hmc_inst.sync_mode_5 = "asynchronous";
defparam hmc_inst.test_mode = "normal_mode";
defparam hmc_inst.thld_jar1_0 = "threshold_32";
defparam hmc_inst.thld_jar1_1 = "threshold_32";
defparam hmc_inst.thld_jar1_2 = "threshold_32";
defparam hmc_inst.thld_jar1_3 = "threshold_32";
defparam hmc_inst.thld_jar1_4 = "threshold_32";
defparam hmc_inst.thld_jar1_5 = "threshold_32";
defparam hmc_inst.thld_jar2_0 = "threshold_16";
defparam hmc_inst.thld_jar2_1 = "threshold_16";
defparam hmc_inst.thld_jar2_2 = "threshold_16";
defparam hmc_inst.thld_jar2_3 = "threshold_16";
defparam hmc_inst.thld_jar2_4 = "threshold_16";
defparam hmc_inst.thld_jar2_5 = "threshold_16";
defparam hmc_inst.use_almost_empty_0 = "empty";
defparam hmc_inst.use_almost_empty_1 = "empty";
defparam hmc_inst.use_almost_empty_2 = "empty";
defparam hmc_inst.use_almost_empty_3 = "empty";
defparam hmc_inst.user_ecc_en = "disable";
defparam hmc_inst.user_priority_0 = "priority_1";
defparam hmc_inst.user_priority_1 = "priority_1";
defparam hmc_inst.user_priority_2 = "priority_1";
defparam hmc_inst.user_priority_3 = "priority_1";
defparam hmc_inst.user_priority_4 = "priority_1";
defparam hmc_inst.user_priority_5 = "priority_1";
defparam hmc_inst.wfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo0_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo1_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo2_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo3_rdy_almost_full = "not_full";
defparam hmc_inst.wr_dwidth_0 = "dwidth_0";
defparam hmc_inst.wr_dwidth_1 = "dwidth_0";
defparam hmc_inst.wr_dwidth_2 = "dwidth_0";
defparam hmc_inst.wr_dwidth_3 = "dwidth_0";
defparam hmc_inst.wr_dwidth_4 = "dwidth_0";
defparam hmc_inst.wr_dwidth_5 = "dwidth_0";
defparam hmc_inst.wr_fifo_in_use_0 = "false";
defparam hmc_inst.wr_fifo_in_use_1 = "false";
defparam hmc_inst.wr_fifo_in_use_2 = "false";
defparam hmc_inst.wr_fifo_in_use_3 = "false";
defparam hmc_inst.wr_port_info_0 = "use_no";
defparam hmc_inst.wr_port_info_1 = "use_no";
defparam hmc_inst.wr_port_info_2 = "use_no";
defparam hmc_inst.wr_port_info_3 = "use_no";
defparam hmc_inst.wr_port_info_4 = "use_no";
defparam hmc_inst.wr_port_info_5 = "use_no";
defparam hmc_inst.write_odt_chip = "write_chip0_odt0_chip1";

endmodule

module system_altera_mem_if_oct_cyclonev (
	parallelterminationcontrol,
	seriesterminationcontrol,
	oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[15:0] parallelterminationcontrol;
output 	[15:0] seriesterminationcontrol;
input 	oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sd1a_0~O_CLKUSRDFTOUT ;
wire \wire_sd1a_serdataout[0] ;

wire [15:0] sd2a_0_PARALLELTERMINATIONCONTROL_bus;
wire [15:0] sd2a_0_SERIESTERMINATIONCONTROL_bus;

assign parallelterminationcontrol[0] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[0];
assign parallelterminationcontrol[1] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[1];
assign parallelterminationcontrol[2] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[2];
assign parallelterminationcontrol[3] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[3];
assign parallelterminationcontrol[4] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[4];
assign parallelterminationcontrol[5] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[5];
assign parallelterminationcontrol[6] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[6];
assign parallelterminationcontrol[7] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[7];
assign parallelterminationcontrol[8] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[8];
assign parallelterminationcontrol[9] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[9];
assign parallelterminationcontrol[10] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[10];
assign parallelterminationcontrol[11] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[11];
assign parallelterminationcontrol[12] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[12];
assign parallelterminationcontrol[13] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[13];
assign parallelterminationcontrol[14] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[14];
assign parallelterminationcontrol[15] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[15];

assign seriesterminationcontrol[0] = sd2a_0_SERIESTERMINATIONCONTROL_bus[0];
assign seriesterminationcontrol[1] = sd2a_0_SERIESTERMINATIONCONTROL_bus[1];
assign seriesterminationcontrol[2] = sd2a_0_SERIESTERMINATIONCONTROL_bus[2];
assign seriesterminationcontrol[3] = sd2a_0_SERIESTERMINATIONCONTROL_bus[3];
assign seriesterminationcontrol[4] = sd2a_0_SERIESTERMINATIONCONTROL_bus[4];
assign seriesterminationcontrol[5] = sd2a_0_SERIESTERMINATIONCONTROL_bus[5];
assign seriesterminationcontrol[6] = sd2a_0_SERIESTERMINATIONCONTROL_bus[6];
assign seriesterminationcontrol[7] = sd2a_0_SERIESTERMINATIONCONTROL_bus[7];
assign seriesterminationcontrol[8] = sd2a_0_SERIESTERMINATIONCONTROL_bus[8];
assign seriesterminationcontrol[9] = sd2a_0_SERIESTERMINATIONCONTROL_bus[9];
assign seriesterminationcontrol[10] = sd2a_0_SERIESTERMINATIONCONTROL_bus[10];
assign seriesterminationcontrol[11] = sd2a_0_SERIESTERMINATIONCONTROL_bus[11];
assign seriesterminationcontrol[12] = sd2a_0_SERIESTERMINATIONCONTROL_bus[12];
assign seriesterminationcontrol[13] = sd2a_0_SERIESTERMINATIONCONTROL_bus[13];
assign seriesterminationcontrol[14] = sd2a_0_SERIESTERMINATIONCONTROL_bus[14];
assign seriesterminationcontrol[15] = sd2a_0_SERIESTERMINATIONCONTROL_bus[15];

cyclonev_termination_logic sd2a_0(
	.s2pload(gnd),
	.scanclk(gnd),
	.scanenable(gnd),
	.serdata(\wire_sd1a_serdataout[0] ),
	.enser(4'b0000),
	.parallelterminationcontrol(sd2a_0_PARALLELTERMINATIONCONTROL_bus),
	.seriesterminationcontrol(sd2a_0_SERIESTERMINATIONCONTROL_bus));

cyclonev_termination sd1a_0(
	.clkenusr(gnd),
	.clkusr(gnd),
	.enserusr(gnd),
	.nclrusr(gnd),
	.rzqin(oct_rzqin),
	.scanclk(gnd),
	.scanen(gnd),
	.scanin(gnd),
	.serdatafromcore(gnd),
	.serdatain(gnd),
	.otherenser(10'b0000000000),
	.clkusrdftout(\sd1a_0~O_CLKUSRDFTOUT ),
	.compoutrdn(),
	.compoutrup(),
	.enserout(),
	.scanout(),
	.serdataout(\wire_sd1a_serdataout[0] ),
	.serdatatocore());

endmodule

module system_hps_sdram_p0 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid_0,
	ctl_reset_n,
	afi_rdata_0,
	afi_rdata_1,
	afi_rdata_2,
	afi_rdata_3,
	afi_rdata_4,
	afi_rdata_5,
	afi_rdata_6,
	afi_rdata_7,
	afi_rdata_8,
	afi_rdata_9,
	afi_rdata_10,
	afi_rdata_11,
	afi_rdata_12,
	afi_rdata_13,
	afi_rdata_14,
	afi_rdata_15,
	afi_rdata_16,
	afi_rdata_17,
	afi_rdata_18,
	afi_rdata_19,
	afi_rdata_20,
	afi_rdata_21,
	afi_rdata_22,
	afi_rdata_23,
	afi_rdata_24,
	afi_rdata_25,
	afi_rdata_26,
	afi_rdata_27,
	afi_rdata_28,
	afi_rdata_29,
	afi_rdata_30,
	afi_rdata_31,
	afi_rdata_32,
	afi_rdata_33,
	afi_rdata_34,
	afi_rdata_35,
	afi_rdata_36,
	afi_rdata_37,
	afi_rdata_38,
	afi_rdata_39,
	afi_rdata_40,
	afi_rdata_41,
	afi_rdata_42,
	afi_rdata_43,
	afi_rdata_44,
	afi_rdata_45,
	afi_rdata_46,
	afi_rdata_47,
	afi_rdata_48,
	afi_rdata_49,
	afi_rdata_50,
	afi_rdata_51,
	afi_rdata_52,
	afi_rdata_53,
	afi_rdata_54,
	afi_rdata_55,
	afi_rdata_56,
	afi_rdata_57,
	afi_rdata_58,
	afi_rdata_59,
	afi_rdata_60,
	afi_rdata_61,
	afi_rdata_62,
	afi_rdata_63,
	afi_rdata_64,
	afi_rdata_65,
	afi_rdata_66,
	afi_rdata_67,
	afi_rdata_68,
	afi_rdata_69,
	afi_rdata_70,
	afi_rdata_71,
	afi_rdata_72,
	afi_rdata_73,
	afi_rdata_74,
	afi_rdata_75,
	afi_rdata_76,
	afi_rdata_77,
	afi_rdata_78,
	afi_rdata_79,
	afi_wlat_0,
	afi_wlat_1,
	afi_wlat_2,
	afi_wlat_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n_0,
	afi_ras_n_0,
	afi_rst_n_0,
	afi_we_n_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_addr_14,
	afi_addr_15,
	afi_addr_16,
	afi_addr_17,
	afi_addr_18,
	afi_addr_19,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_cke_0,
	afi_cke_1,
	afi_cs_n_0,
	afi_cs_n_1,
	afi_dm_int_0,
	afi_dm_int_1,
	afi_dm_int_2,
	afi_dm_int_3,
	afi_dm_int_4,
	afi_dm_int_5,
	afi_dm_int_6,
	afi_dm_int_7,
	afi_dm_int_8,
	afi_dm_int_9,
	afi_dqs_burst_0,
	afi_dqs_burst_1,
	afi_dqs_burst_2,
	afi_dqs_burst_3,
	afi_dqs_burst_4,
	afi_odt_0,
	afi_odt_1,
	afi_rdata_en_0,
	afi_rdata_en_1,
	afi_rdata_en_2,
	afi_rdata_en_3,
	afi_rdata_en_4,
	afi_rdata_en_full_0,
	afi_rdata_en_full_1,
	afi_rdata_en_full_2,
	afi_rdata_en_full_3,
	afi_rdata_en_full_4,
	afi_wdata_int_0,
	afi_wdata_int_1,
	afi_wdata_int_2,
	afi_wdata_int_3,
	afi_wdata_int_4,
	afi_wdata_int_5,
	afi_wdata_int_6,
	afi_wdata_int_7,
	afi_wdata_int_8,
	afi_wdata_int_9,
	afi_wdata_int_10,
	afi_wdata_int_11,
	afi_wdata_int_12,
	afi_wdata_int_13,
	afi_wdata_int_14,
	afi_wdata_int_15,
	afi_wdata_int_16,
	afi_wdata_int_17,
	afi_wdata_int_18,
	afi_wdata_int_19,
	afi_wdata_int_20,
	afi_wdata_int_21,
	afi_wdata_int_22,
	afi_wdata_int_23,
	afi_wdata_int_24,
	afi_wdata_int_25,
	afi_wdata_int_26,
	afi_wdata_int_27,
	afi_wdata_int_28,
	afi_wdata_int_29,
	afi_wdata_int_30,
	afi_wdata_int_31,
	afi_wdata_int_32,
	afi_wdata_int_33,
	afi_wdata_int_34,
	afi_wdata_int_35,
	afi_wdata_int_36,
	afi_wdata_int_37,
	afi_wdata_int_38,
	afi_wdata_int_39,
	afi_wdata_int_40,
	afi_wdata_int_41,
	afi_wdata_int_42,
	afi_wdata_int_43,
	afi_wdata_int_44,
	afi_wdata_int_45,
	afi_wdata_int_46,
	afi_wdata_int_47,
	afi_wdata_int_48,
	afi_wdata_int_49,
	afi_wdata_int_50,
	afi_wdata_int_51,
	afi_wdata_int_52,
	afi_wdata_int_53,
	afi_wdata_int_54,
	afi_wdata_int_55,
	afi_wdata_int_56,
	afi_wdata_int_57,
	afi_wdata_int_58,
	afi_wdata_int_59,
	afi_wdata_int_60,
	afi_wdata_int_61,
	afi_wdata_int_62,
	afi_wdata_int_63,
	afi_wdata_int_64,
	afi_wdata_int_65,
	afi_wdata_int_66,
	afi_wdata_int_67,
	afi_wdata_int_68,
	afi_wdata_int_69,
	afi_wdata_int_70,
	afi_wdata_int_71,
	afi_wdata_int_72,
	afi_wdata_int_73,
	afi_wdata_int_74,
	afi_wdata_int_75,
	afi_wdata_int_76,
	afi_wdata_int_77,
	afi_wdata_int_78,
	afi_wdata_int_79,
	afi_wdata_valid_0,
	afi_wdata_valid_1,
	afi_wdata_valid_2,
	afi_wdata_valid_3,
	afi_wdata_valid_4,
	cfg_addlat_wire_0,
	cfg_addlat_wire_1,
	cfg_addlat_wire_2,
	cfg_addlat_wire_3,
	cfg_addlat_wire_4,
	cfg_bankaddrwidth_wire_0,
	cfg_bankaddrwidth_wire_1,
	cfg_bankaddrwidth_wire_2,
	cfg_caswrlat_wire_0,
	cfg_caswrlat_wire_1,
	cfg_caswrlat_wire_2,
	cfg_caswrlat_wire_3,
	cfg_coladdrwidth_wire_0,
	cfg_coladdrwidth_wire_1,
	cfg_coladdrwidth_wire_2,
	cfg_coladdrwidth_wire_3,
	cfg_coladdrwidth_wire_4,
	cfg_csaddrwidth_wire_0,
	cfg_csaddrwidth_wire_1,
	cfg_csaddrwidth_wire_2,
	cfg_devicewidth_wire_0,
	cfg_devicewidth_wire_1,
	cfg_devicewidth_wire_2,
	cfg_devicewidth_wire_3,
	cfg_interfacewidth_wire_0,
	cfg_interfacewidth_wire_1,
	cfg_interfacewidth_wire_2,
	cfg_interfacewidth_wire_3,
	cfg_interfacewidth_wire_4,
	cfg_interfacewidth_wire_5,
	cfg_interfacewidth_wire_6,
	cfg_interfacewidth_wire_7,
	cfg_rowaddrwidth_wire_0,
	cfg_rowaddrwidth_wire_1,
	cfg_rowaddrwidth_wire_2,
	cfg_rowaddrwidth_wire_3,
	cfg_rowaddrwidth_wire_4,
	cfg_tcl_wire_0,
	cfg_tcl_wire_1,
	cfg_tcl_wire_2,
	cfg_tcl_wire_3,
	cfg_tcl_wire_4,
	cfg_tmrd_wire_0,
	cfg_tmrd_wire_1,
	cfg_tmrd_wire_2,
	cfg_tmrd_wire_3,
	cfg_trefi_wire_0,
	cfg_trefi_wire_1,
	cfg_trefi_wire_2,
	cfg_trefi_wire_3,
	cfg_trefi_wire_4,
	cfg_trefi_wire_5,
	cfg_trefi_wire_6,
	cfg_trefi_wire_7,
	cfg_trefi_wire_8,
	cfg_trefi_wire_9,
	cfg_trefi_wire_10,
	cfg_trefi_wire_11,
	cfg_trefi_wire_12,
	cfg_trfc_wire_0,
	cfg_trfc_wire_1,
	cfg_trfc_wire_2,
	cfg_trfc_wire_3,
	cfg_trfc_wire_4,
	cfg_trfc_wire_5,
	cfg_trfc_wire_6,
	cfg_trfc_wire_7,
	cfg_twr_wire_0,
	cfg_twr_wire_1,
	cfg_twr_wire_2,
	cfg_twr_wire_3,
	afi_mem_clk_disable_0,
	cfg_dramconfig_wire_0,
	cfg_dramconfig_wire_1,
	cfg_dramconfig_wire_2,
	cfg_dramconfig_wire_3,
	cfg_dramconfig_wire_4,
	cfg_dramconfig_wire_5,
	cfg_dramconfig_wire_6,
	cfg_dramconfig_wire_7,
	cfg_dramconfig_wire_8,
	cfg_dramconfig_wire_9,
	cfg_dramconfig_wire_10,
	cfg_dramconfig_wire_11,
	cfg_dramconfig_wire_12,
	cfg_dramconfig_wire_13,
	cfg_dramconfig_wire_14,
	cfg_dramconfig_wire_15,
	cfg_dramconfig_wire_16,
	cfg_dramconfig_wire_17,
	cfg_dramconfig_wire_18,
	cfg_dramconfig_wire_19,
	cfg_dramconfig_wire_20,
	leveled_dqs_clocks_0,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	afi_rdata_valid_0;
output 	ctl_reset_n;
output 	afi_rdata_0;
output 	afi_rdata_1;
output 	afi_rdata_2;
output 	afi_rdata_3;
output 	afi_rdata_4;
output 	afi_rdata_5;
output 	afi_rdata_6;
output 	afi_rdata_7;
output 	afi_rdata_8;
output 	afi_rdata_9;
output 	afi_rdata_10;
output 	afi_rdata_11;
output 	afi_rdata_12;
output 	afi_rdata_13;
output 	afi_rdata_14;
output 	afi_rdata_15;
output 	afi_rdata_16;
output 	afi_rdata_17;
output 	afi_rdata_18;
output 	afi_rdata_19;
output 	afi_rdata_20;
output 	afi_rdata_21;
output 	afi_rdata_22;
output 	afi_rdata_23;
output 	afi_rdata_24;
output 	afi_rdata_25;
output 	afi_rdata_26;
output 	afi_rdata_27;
output 	afi_rdata_28;
output 	afi_rdata_29;
output 	afi_rdata_30;
output 	afi_rdata_31;
output 	afi_rdata_32;
output 	afi_rdata_33;
output 	afi_rdata_34;
output 	afi_rdata_35;
output 	afi_rdata_36;
output 	afi_rdata_37;
output 	afi_rdata_38;
output 	afi_rdata_39;
output 	afi_rdata_40;
output 	afi_rdata_41;
output 	afi_rdata_42;
output 	afi_rdata_43;
output 	afi_rdata_44;
output 	afi_rdata_45;
output 	afi_rdata_46;
output 	afi_rdata_47;
output 	afi_rdata_48;
output 	afi_rdata_49;
output 	afi_rdata_50;
output 	afi_rdata_51;
output 	afi_rdata_52;
output 	afi_rdata_53;
output 	afi_rdata_54;
output 	afi_rdata_55;
output 	afi_rdata_56;
output 	afi_rdata_57;
output 	afi_rdata_58;
output 	afi_rdata_59;
output 	afi_rdata_60;
output 	afi_rdata_61;
output 	afi_rdata_62;
output 	afi_rdata_63;
output 	afi_rdata_64;
output 	afi_rdata_65;
output 	afi_rdata_66;
output 	afi_rdata_67;
output 	afi_rdata_68;
output 	afi_rdata_69;
output 	afi_rdata_70;
output 	afi_rdata_71;
output 	afi_rdata_72;
output 	afi_rdata_73;
output 	afi_rdata_74;
output 	afi_rdata_75;
output 	afi_rdata_76;
output 	afi_rdata_77;
output 	afi_rdata_78;
output 	afi_rdata_79;
output 	afi_wlat_0;
output 	afi_wlat_1;
output 	afi_wlat_2;
output 	afi_wlat_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	afi_cas_n_0;
input 	afi_ras_n_0;
input 	afi_rst_n_0;
input 	afi_we_n_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_addr_14;
input 	afi_addr_15;
input 	afi_addr_16;
input 	afi_addr_17;
input 	afi_addr_18;
input 	afi_addr_19;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_cke_0;
input 	afi_cke_1;
input 	afi_cs_n_0;
input 	afi_cs_n_1;
input 	afi_dm_int_0;
input 	afi_dm_int_1;
input 	afi_dm_int_2;
input 	afi_dm_int_3;
input 	afi_dm_int_4;
input 	afi_dm_int_5;
input 	afi_dm_int_6;
input 	afi_dm_int_7;
input 	afi_dm_int_8;
input 	afi_dm_int_9;
input 	afi_dqs_burst_0;
input 	afi_dqs_burst_1;
input 	afi_dqs_burst_2;
input 	afi_dqs_burst_3;
input 	afi_dqs_burst_4;
input 	afi_odt_0;
input 	afi_odt_1;
input 	afi_rdata_en_0;
input 	afi_rdata_en_1;
input 	afi_rdata_en_2;
input 	afi_rdata_en_3;
input 	afi_rdata_en_4;
input 	afi_rdata_en_full_0;
input 	afi_rdata_en_full_1;
input 	afi_rdata_en_full_2;
input 	afi_rdata_en_full_3;
input 	afi_rdata_en_full_4;
input 	afi_wdata_int_0;
input 	afi_wdata_int_1;
input 	afi_wdata_int_2;
input 	afi_wdata_int_3;
input 	afi_wdata_int_4;
input 	afi_wdata_int_5;
input 	afi_wdata_int_6;
input 	afi_wdata_int_7;
input 	afi_wdata_int_8;
input 	afi_wdata_int_9;
input 	afi_wdata_int_10;
input 	afi_wdata_int_11;
input 	afi_wdata_int_12;
input 	afi_wdata_int_13;
input 	afi_wdata_int_14;
input 	afi_wdata_int_15;
input 	afi_wdata_int_16;
input 	afi_wdata_int_17;
input 	afi_wdata_int_18;
input 	afi_wdata_int_19;
input 	afi_wdata_int_20;
input 	afi_wdata_int_21;
input 	afi_wdata_int_22;
input 	afi_wdata_int_23;
input 	afi_wdata_int_24;
input 	afi_wdata_int_25;
input 	afi_wdata_int_26;
input 	afi_wdata_int_27;
input 	afi_wdata_int_28;
input 	afi_wdata_int_29;
input 	afi_wdata_int_30;
input 	afi_wdata_int_31;
input 	afi_wdata_int_32;
input 	afi_wdata_int_33;
input 	afi_wdata_int_34;
input 	afi_wdata_int_35;
input 	afi_wdata_int_36;
input 	afi_wdata_int_37;
input 	afi_wdata_int_38;
input 	afi_wdata_int_39;
input 	afi_wdata_int_40;
input 	afi_wdata_int_41;
input 	afi_wdata_int_42;
input 	afi_wdata_int_43;
input 	afi_wdata_int_44;
input 	afi_wdata_int_45;
input 	afi_wdata_int_46;
input 	afi_wdata_int_47;
input 	afi_wdata_int_48;
input 	afi_wdata_int_49;
input 	afi_wdata_int_50;
input 	afi_wdata_int_51;
input 	afi_wdata_int_52;
input 	afi_wdata_int_53;
input 	afi_wdata_int_54;
input 	afi_wdata_int_55;
input 	afi_wdata_int_56;
input 	afi_wdata_int_57;
input 	afi_wdata_int_58;
input 	afi_wdata_int_59;
input 	afi_wdata_int_60;
input 	afi_wdata_int_61;
input 	afi_wdata_int_62;
input 	afi_wdata_int_63;
input 	afi_wdata_int_64;
input 	afi_wdata_int_65;
input 	afi_wdata_int_66;
input 	afi_wdata_int_67;
input 	afi_wdata_int_68;
input 	afi_wdata_int_69;
input 	afi_wdata_int_70;
input 	afi_wdata_int_71;
input 	afi_wdata_int_72;
input 	afi_wdata_int_73;
input 	afi_wdata_int_74;
input 	afi_wdata_int_75;
input 	afi_wdata_int_76;
input 	afi_wdata_int_77;
input 	afi_wdata_int_78;
input 	afi_wdata_int_79;
input 	afi_wdata_valid_0;
input 	afi_wdata_valid_1;
input 	afi_wdata_valid_2;
input 	afi_wdata_valid_3;
input 	afi_wdata_valid_4;
input 	cfg_addlat_wire_0;
input 	cfg_addlat_wire_1;
input 	cfg_addlat_wire_2;
input 	cfg_addlat_wire_3;
input 	cfg_addlat_wire_4;
input 	cfg_bankaddrwidth_wire_0;
input 	cfg_bankaddrwidth_wire_1;
input 	cfg_bankaddrwidth_wire_2;
input 	cfg_caswrlat_wire_0;
input 	cfg_caswrlat_wire_1;
input 	cfg_caswrlat_wire_2;
input 	cfg_caswrlat_wire_3;
input 	cfg_coladdrwidth_wire_0;
input 	cfg_coladdrwidth_wire_1;
input 	cfg_coladdrwidth_wire_2;
input 	cfg_coladdrwidth_wire_3;
input 	cfg_coladdrwidth_wire_4;
input 	cfg_csaddrwidth_wire_0;
input 	cfg_csaddrwidth_wire_1;
input 	cfg_csaddrwidth_wire_2;
input 	cfg_devicewidth_wire_0;
input 	cfg_devicewidth_wire_1;
input 	cfg_devicewidth_wire_2;
input 	cfg_devicewidth_wire_3;
input 	cfg_interfacewidth_wire_0;
input 	cfg_interfacewidth_wire_1;
input 	cfg_interfacewidth_wire_2;
input 	cfg_interfacewidth_wire_3;
input 	cfg_interfacewidth_wire_4;
input 	cfg_interfacewidth_wire_5;
input 	cfg_interfacewidth_wire_6;
input 	cfg_interfacewidth_wire_7;
input 	cfg_rowaddrwidth_wire_0;
input 	cfg_rowaddrwidth_wire_1;
input 	cfg_rowaddrwidth_wire_2;
input 	cfg_rowaddrwidth_wire_3;
input 	cfg_rowaddrwidth_wire_4;
input 	cfg_tcl_wire_0;
input 	cfg_tcl_wire_1;
input 	cfg_tcl_wire_2;
input 	cfg_tcl_wire_3;
input 	cfg_tcl_wire_4;
input 	cfg_tmrd_wire_0;
input 	cfg_tmrd_wire_1;
input 	cfg_tmrd_wire_2;
input 	cfg_tmrd_wire_3;
input 	cfg_trefi_wire_0;
input 	cfg_trefi_wire_1;
input 	cfg_trefi_wire_2;
input 	cfg_trefi_wire_3;
input 	cfg_trefi_wire_4;
input 	cfg_trefi_wire_5;
input 	cfg_trefi_wire_6;
input 	cfg_trefi_wire_7;
input 	cfg_trefi_wire_8;
input 	cfg_trefi_wire_9;
input 	cfg_trefi_wire_10;
input 	cfg_trefi_wire_11;
input 	cfg_trefi_wire_12;
input 	cfg_trfc_wire_0;
input 	cfg_trfc_wire_1;
input 	cfg_trfc_wire_2;
input 	cfg_trfc_wire_3;
input 	cfg_trfc_wire_4;
input 	cfg_trfc_wire_5;
input 	cfg_trfc_wire_6;
input 	cfg_trfc_wire_7;
input 	cfg_twr_wire_0;
input 	cfg_twr_wire_1;
input 	cfg_twr_wire_2;
input 	cfg_twr_wire_3;
input 	afi_mem_clk_disable_0;
input 	cfg_dramconfig_wire_0;
input 	cfg_dramconfig_wire_1;
input 	cfg_dramconfig_wire_2;
input 	cfg_dramconfig_wire_3;
input 	cfg_dramconfig_wire_4;
input 	cfg_dramconfig_wire_5;
input 	cfg_dramconfig_wire_6;
input 	cfg_dramconfig_wire_7;
input 	cfg_dramconfig_wire_8;
input 	cfg_dramconfig_wire_9;
input 	cfg_dramconfig_wire_10;
input 	cfg_dramconfig_wire_11;
input 	cfg_dramconfig_wire_12;
input 	cfg_dramconfig_wire_13;
input 	cfg_dramconfig_wire_14;
input 	cfg_dramconfig_wire_15;
input 	cfg_dramconfig_wire_16;
input 	cfg_dramconfig_wire_17;
input 	cfg_dramconfig_wire_18;
input 	cfg_dramconfig_wire_19;
input 	cfg_dramconfig_wire_20;
output 	leveled_dqs_clocks_0;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_hps_sdram_p0_acv_hard_memphy umemphy(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(afi_cal_fail),
	.afi_cal_success(afi_cal_success),
	.afi_rdata_valid({afi_rdata_valid_0}),
	.ctl_reset_n(ctl_reset_n),
	.afi_rdata({afi_rdata_79,afi_rdata_78,afi_rdata_77,afi_rdata_76,afi_rdata_75,afi_rdata_74,afi_rdata_73,afi_rdata_72,afi_rdata_71,afi_rdata_70,afi_rdata_69,afi_rdata_68,afi_rdata_67,afi_rdata_66,afi_rdata_65,afi_rdata_64,afi_rdata_63,afi_rdata_62,afi_rdata_61,afi_rdata_60,afi_rdata_59,
afi_rdata_58,afi_rdata_57,afi_rdata_56,afi_rdata_55,afi_rdata_54,afi_rdata_53,afi_rdata_52,afi_rdata_51,afi_rdata_50,afi_rdata_49,afi_rdata_48,afi_rdata_47,afi_rdata_46,afi_rdata_45,afi_rdata_44,afi_rdata_43,afi_rdata_42,afi_rdata_41,afi_rdata_40,afi_rdata_39,afi_rdata_38,
afi_rdata_37,afi_rdata_36,afi_rdata_35,afi_rdata_34,afi_rdata_33,afi_rdata_32,afi_rdata_31,afi_rdata_30,afi_rdata_29,afi_rdata_28,afi_rdata_27,afi_rdata_26,afi_rdata_25,afi_rdata_24,afi_rdata_23,afi_rdata_22,afi_rdata_21,afi_rdata_20,afi_rdata_19,afi_rdata_18,afi_rdata_17,
afi_rdata_16,afi_rdata_15,afi_rdata_14,afi_rdata_13,afi_rdata_12,afi_rdata_11,afi_rdata_10,afi_rdata_9,afi_rdata_8,afi_rdata_7,afi_rdata_6,afi_rdata_5,afi_rdata_4,afi_rdata_3,afi_rdata_2,afi_rdata_1,afi_rdata_0}),
	.afi_wlat({afi_wlat_3,afi_wlat_2,afi_wlat_1,afi_wlat_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n({afi_cas_n_0}),
	.afi_ras_n({afi_ras_n_0}),
	.afi_rst_n({afi_rst_n_0}),
	.afi_we_n({afi_we_n_0}),
	.afi_addr({afi_addr_19,afi_addr_18,afi_addr_17,afi_addr_16,afi_addr_15,afi_addr_14,afi_addr_13,afi_addr_12,afi_addr_11,afi_addr_10,afi_addr_9,afi_addr_8,afi_addr_7,afi_addr_6,afi_addr_5,afi_addr_4,afi_addr_3,afi_addr_2,afi_addr_1,afi_addr_0}),
	.afi_ba({afi_ba_2,afi_ba_1,afi_ba_0}),
	.afi_cke({afi_cke_1,afi_cke_0}),
	.afi_cs_n({afi_cs_n_1,afi_cs_n_0}),
	.afi_dm({afi_dm_int_9,afi_dm_int_8,afi_dm_int_7,afi_dm_int_6,afi_dm_int_5,afi_dm_int_4,afi_dm_int_3,afi_dm_int_2,afi_dm_int_1,afi_dm_int_0}),
	.afi_dqs_burst({afi_dqs_burst_4,afi_dqs_burst_3,afi_dqs_burst_2,afi_dqs_burst_1,afi_dqs_burst_0}),
	.afi_odt({afi_odt_1,afi_odt_0}),
	.afi_rdata_en({afi_rdata_en_4,afi_rdata_en_3,afi_rdata_en_2,afi_rdata_en_1,afi_rdata_en_0}),
	.afi_rdata_en_full({afi_rdata_en_full_4,afi_rdata_en_full_3,afi_rdata_en_full_2,afi_rdata_en_full_1,afi_rdata_en_full_0}),
	.afi_wdata({afi_wdata_int_79,afi_wdata_int_78,afi_wdata_int_77,afi_wdata_int_76,afi_wdata_int_75,afi_wdata_int_74,afi_wdata_int_73,afi_wdata_int_72,afi_wdata_int_71,afi_wdata_int_70,afi_wdata_int_69,afi_wdata_int_68,afi_wdata_int_67,afi_wdata_int_66,afi_wdata_int_65,afi_wdata_int_64,
afi_wdata_int_63,afi_wdata_int_62,afi_wdata_int_61,afi_wdata_int_60,afi_wdata_int_59,afi_wdata_int_58,afi_wdata_int_57,afi_wdata_int_56,afi_wdata_int_55,afi_wdata_int_54,afi_wdata_int_53,afi_wdata_int_52,afi_wdata_int_51,afi_wdata_int_50,afi_wdata_int_49,afi_wdata_int_48,
afi_wdata_int_47,afi_wdata_int_46,afi_wdata_int_45,afi_wdata_int_44,afi_wdata_int_43,afi_wdata_int_42,afi_wdata_int_41,afi_wdata_int_40,afi_wdata_int_39,afi_wdata_int_38,afi_wdata_int_37,afi_wdata_int_36,afi_wdata_int_35,afi_wdata_int_34,afi_wdata_int_33,afi_wdata_int_32,
afi_wdata_int_31,afi_wdata_int_30,afi_wdata_int_29,afi_wdata_int_28,afi_wdata_int_27,afi_wdata_int_26,afi_wdata_int_25,afi_wdata_int_24,afi_wdata_int_23,afi_wdata_int_22,afi_wdata_int_21,afi_wdata_int_20,afi_wdata_int_19,afi_wdata_int_18,afi_wdata_int_17,afi_wdata_int_16,
afi_wdata_int_15,afi_wdata_int_14,afi_wdata_int_13,afi_wdata_int_12,afi_wdata_int_11,afi_wdata_int_10,afi_wdata_int_9,afi_wdata_int_8,afi_wdata_int_7,afi_wdata_int_6,afi_wdata_int_5,afi_wdata_int_4,afi_wdata_int_3,afi_wdata_int_2,afi_wdata_int_1,afi_wdata_int_0}),
	.afi_wdata_valid({afi_wdata_valid_4,afi_wdata_valid_3,afi_wdata_valid_2,afi_wdata_valid_1,afi_wdata_valid_0}),
	.cfg_addlat({gnd,gnd,gnd,cfg_addlat_wire_4,cfg_addlat_wire_3,cfg_addlat_wire_2,cfg_addlat_wire_1,cfg_addlat_wire_0}),
	.cfg_bankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth_wire_2,cfg_bankaddrwidth_wire_1,cfg_bankaddrwidth_wire_0}),
	.cfg_caswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat_wire_3,cfg_caswrlat_wire_2,cfg_caswrlat_wire_1,cfg_caswrlat_wire_0}),
	.cfg_coladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth_wire_4,cfg_coladdrwidth_wire_3,cfg_coladdrwidth_wire_2,cfg_coladdrwidth_wire_1,cfg_coladdrwidth_wire_0}),
	.cfg_csaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth_wire_2,cfg_csaddrwidth_wire_1,cfg_csaddrwidth_wire_0}),
	.cfg_devicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth_wire_3,cfg_devicewidth_wire_2,cfg_devicewidth_wire_1,cfg_devicewidth_wire_0}),
	.cfg_interfacewidth({cfg_interfacewidth_wire_7,cfg_interfacewidth_wire_6,cfg_interfacewidth_wire_5,cfg_interfacewidth_wire_4,cfg_interfacewidth_wire_3,cfg_interfacewidth_wire_2,cfg_interfacewidth_wire_1,cfg_interfacewidth_wire_0}),
	.cfg_rowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth_wire_4,cfg_rowaddrwidth_wire_3,cfg_rowaddrwidth_wire_2,cfg_rowaddrwidth_wire_1,cfg_rowaddrwidth_wire_0}),
	.cfg_tcl({gnd,gnd,gnd,cfg_tcl_wire_4,cfg_tcl_wire_3,cfg_tcl_wire_2,cfg_tcl_wire_1,cfg_tcl_wire_0}),
	.cfg_tmrd({gnd,gnd,gnd,gnd,cfg_tmrd_wire_3,cfg_tmrd_wire_2,cfg_tmrd_wire_1,cfg_tmrd_wire_0}),
	.cfg_trefi({gnd,gnd,gnd,cfg_trefi_wire_12,cfg_trefi_wire_11,cfg_trefi_wire_10,cfg_trefi_wire_9,cfg_trefi_wire_8,cfg_trefi_wire_7,cfg_trefi_wire_6,cfg_trefi_wire_5,cfg_trefi_wire_4,cfg_trefi_wire_3,cfg_trefi_wire_2,cfg_trefi_wire_1,cfg_trefi_wire_0}),
	.cfg_trfc({cfg_trfc_wire_7,cfg_trfc_wire_6,cfg_trfc_wire_5,cfg_trfc_wire_4,cfg_trfc_wire_3,cfg_trfc_wire_2,cfg_trfc_wire_1,cfg_trfc_wire_0}),
	.cfg_twr({gnd,gnd,gnd,gnd,cfg_twr_wire_3,cfg_twr_wire_2,cfg_twr_wire_1,cfg_twr_wire_0}),
	.afi_mem_clk_disable({afi_mem_clk_disable_0}),
	.cfg_dramconfig({gnd,gnd,gnd,cfg_dramconfig_wire_20,cfg_dramconfig_wire_19,cfg_dramconfig_wire_18,cfg_dramconfig_wire_17,cfg_dramconfig_wire_16,cfg_dramconfig_wire_15,cfg_dramconfig_wire_14,cfg_dramconfig_wire_13,cfg_dramconfig_wire_12,cfg_dramconfig_wire_11,cfg_dramconfig_wire_10,
cfg_dramconfig_wire_9,cfg_dramconfig_wire_8,cfg_dramconfig_wire_7,cfg_dramconfig_wire_6,cfg_dramconfig_wire_5,cfg_dramconfig_wire_4,cfg_dramconfig_wire_3,cfg_dramconfig_wire_2,cfg_dramconfig_wire_1,cfg_dramconfig_wire_0}),
	.leveled_dqs_clocks_0(leveled_dqs_clocks_0),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module system_hps_sdram_p0_acv_hard_memphy (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	leveled_dqs_clocks_0,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	[0:0] afi_rdata_valid;
output 	ctl_reset_n;
output 	[79:0] afi_rdata;
output 	[3:0] afi_wlat;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	[0:0] afi_cas_n;
input 	[0:0] afi_ras_n;
input 	[0:0] afi_rst_n;
input 	[0:0] afi_we_n;
input 	[19:0] afi_addr;
input 	[2:0] afi_ba;
input 	[1:0] afi_cke;
input 	[1:0] afi_cs_n;
input 	[9:0] afi_dm;
input 	[4:0] afi_dqs_burst;
input 	[1:0] afi_odt;
input 	[4:0] afi_rdata_en;
input 	[4:0] afi_rdata_en_full;
input 	[79:0] afi_wdata;
input 	[4:0] afi_wdata_valid;
input 	[7:0] cfg_addlat;
input 	[7:0] cfg_bankaddrwidth;
input 	[7:0] cfg_caswrlat;
input 	[7:0] cfg_coladdrwidth;
input 	[7:0] cfg_csaddrwidth;
input 	[7:0] cfg_devicewidth;
input 	[7:0] cfg_interfacewidth;
input 	[7:0] cfg_rowaddrwidth;
input 	[7:0] cfg_tcl;
input 	[7:0] cfg_tmrd;
input 	[15:0] cfg_trefi;
input 	[7:0] cfg_trfc;
input 	[7:0] cfg_twr;
input 	[0:0] afi_mem_clk_disable;
input 	[23:0] cfg_dramconfig;
output 	leveled_dqs_clocks_0;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \memphy_ldc|leveled_hr_clocks[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \phy_ddio_address[0] ;
wire \phy_ddio_address[1] ;
wire \phy_ddio_address[2] ;
wire \phy_ddio_address[3] ;
wire \phy_ddio_address[4] ;
wire \phy_ddio_address[5] ;
wire \phy_ddio_address[6] ;
wire \phy_ddio_address[7] ;
wire \phy_ddio_address[8] ;
wire \phy_ddio_address[9] ;
wire \phy_ddio_address[10] ;
wire \phy_ddio_address[11] ;
wire \phy_ddio_address[12] ;
wire \phy_ddio_address[13] ;
wire \phy_ddio_address[14] ;
wire \phy_ddio_address[15] ;
wire \phy_ddio_address[16] ;
wire \phy_ddio_address[17] ;
wire \phy_ddio_address[18] ;
wire \phy_ddio_address[19] ;
wire \phy_ddio_address[20] ;
wire \phy_ddio_address[21] ;
wire \phy_ddio_address[22] ;
wire \phy_ddio_address[23] ;
wire \phy_ddio_address[24] ;
wire \phy_ddio_address[25] ;
wire \phy_ddio_address[26] ;
wire \phy_ddio_address[27] ;
wire \phy_ddio_address[28] ;
wire \phy_ddio_address[29] ;
wire \phy_ddio_address[30] ;
wire \phy_ddio_address[31] ;
wire \phy_ddio_address[32] ;
wire \phy_ddio_address[33] ;
wire \phy_ddio_address[34] ;
wire \phy_ddio_address[35] ;
wire \phy_ddio_address[36] ;
wire \phy_ddio_address[37] ;
wire \phy_ddio_address[38] ;
wire \phy_ddio_address[39] ;
wire \phy_ddio_address[40] ;
wire \phy_ddio_address[41] ;
wire \phy_ddio_address[42] ;
wire \phy_ddio_address[43] ;
wire \phy_ddio_address[44] ;
wire \phy_ddio_address[45] ;
wire \phy_ddio_address[46] ;
wire \phy_ddio_address[47] ;
wire \phy_ddio_address[48] ;
wire \phy_ddio_address[49] ;
wire \phy_ddio_address[50] ;
wire \phy_ddio_address[51] ;
wire \phy_ddio_address[52] ;
wire \phy_ddio_address[53] ;
wire \phy_ddio_address[54] ;
wire \phy_ddio_address[55] ;
wire \phy_ddio_address[56] ;
wire \phy_ddio_address[57] ;
wire \phy_ddio_address[58] ;
wire \phy_ddio_address[59] ;
wire \phy_ddio_bank[0] ;
wire \phy_ddio_bank[1] ;
wire \phy_ddio_bank[2] ;
wire \phy_ddio_bank[3] ;
wire \phy_ddio_bank[4] ;
wire \phy_ddio_bank[5] ;
wire \phy_ddio_bank[6] ;
wire \phy_ddio_bank[7] ;
wire \phy_ddio_bank[8] ;
wire \phy_ddio_bank[9] ;
wire \phy_ddio_bank[10] ;
wire \phy_ddio_bank[11] ;
wire \phy_ddio_cas_n[0] ;
wire \phy_ddio_cas_n[1] ;
wire \phy_ddio_cas_n[2] ;
wire \phy_ddio_cas_n[3] ;
wire \phy_ddio_ck[0] ;
wire \phy_ddio_ck[1] ;
wire \phy_ddio_cke[0] ;
wire \phy_ddio_cke[1] ;
wire \phy_ddio_cke[2] ;
wire \phy_ddio_cke[3] ;
wire \phy_ddio_cs_n[0] ;
wire \phy_ddio_cs_n[1] ;
wire \phy_ddio_cs_n[2] ;
wire \phy_ddio_cs_n[3] ;
wire \phy_ddio_dmdout[0] ;
wire \phy_ddio_dmdout[1] ;
wire \phy_ddio_dmdout[2] ;
wire \phy_ddio_dmdout[3] ;
wire \phy_ddio_dmdout[4] ;
wire \phy_ddio_dmdout[5] ;
wire \phy_ddio_dmdout[6] ;
wire \phy_ddio_dmdout[7] ;
wire \phy_ddio_dmdout[8] ;
wire \phy_ddio_dmdout[9] ;
wire \phy_ddio_dmdout[10] ;
wire \phy_ddio_dmdout[11] ;
wire \phy_ddio_dmdout[12] ;
wire \phy_ddio_dmdout[13] ;
wire \phy_ddio_dmdout[14] ;
wire \phy_ddio_dmdout[15] ;
wire \phy_ddio_dqdout[0] ;
wire \phy_ddio_dqdout[1] ;
wire \phy_ddio_dqdout[2] ;
wire \phy_ddio_dqdout[3] ;
wire \phy_ddio_dqdout[4] ;
wire \phy_ddio_dqdout[5] ;
wire \phy_ddio_dqdout[6] ;
wire \phy_ddio_dqdout[7] ;
wire \phy_ddio_dqdout[8] ;
wire \phy_ddio_dqdout[9] ;
wire \phy_ddio_dqdout[10] ;
wire \phy_ddio_dqdout[11] ;
wire \phy_ddio_dqdout[12] ;
wire \phy_ddio_dqdout[13] ;
wire \phy_ddio_dqdout[14] ;
wire \phy_ddio_dqdout[15] ;
wire \phy_ddio_dqdout[16] ;
wire \phy_ddio_dqdout[17] ;
wire \phy_ddio_dqdout[18] ;
wire \phy_ddio_dqdout[19] ;
wire \phy_ddio_dqdout[20] ;
wire \phy_ddio_dqdout[21] ;
wire \phy_ddio_dqdout[22] ;
wire \phy_ddio_dqdout[23] ;
wire \phy_ddio_dqdout[24] ;
wire \phy_ddio_dqdout[25] ;
wire \phy_ddio_dqdout[26] ;
wire \phy_ddio_dqdout[27] ;
wire \phy_ddio_dqdout[28] ;
wire \phy_ddio_dqdout[29] ;
wire \phy_ddio_dqdout[30] ;
wire \phy_ddio_dqdout[31] ;
wire \phy_ddio_dqdout[36] ;
wire \phy_ddio_dqdout[37] ;
wire \phy_ddio_dqdout[38] ;
wire \phy_ddio_dqdout[39] ;
wire \phy_ddio_dqdout[40] ;
wire \phy_ddio_dqdout[41] ;
wire \phy_ddio_dqdout[42] ;
wire \phy_ddio_dqdout[43] ;
wire \phy_ddio_dqdout[44] ;
wire \phy_ddio_dqdout[45] ;
wire \phy_ddio_dqdout[46] ;
wire \phy_ddio_dqdout[47] ;
wire \phy_ddio_dqdout[48] ;
wire \phy_ddio_dqdout[49] ;
wire \phy_ddio_dqdout[50] ;
wire \phy_ddio_dqdout[51] ;
wire \phy_ddio_dqdout[52] ;
wire \phy_ddio_dqdout[53] ;
wire \phy_ddio_dqdout[54] ;
wire \phy_ddio_dqdout[55] ;
wire \phy_ddio_dqdout[56] ;
wire \phy_ddio_dqdout[57] ;
wire \phy_ddio_dqdout[58] ;
wire \phy_ddio_dqdout[59] ;
wire \phy_ddio_dqdout[60] ;
wire \phy_ddio_dqdout[61] ;
wire \phy_ddio_dqdout[62] ;
wire \phy_ddio_dqdout[63] ;
wire \phy_ddio_dqdout[64] ;
wire \phy_ddio_dqdout[65] ;
wire \phy_ddio_dqdout[66] ;
wire \phy_ddio_dqdout[67] ;
wire \phy_ddio_dqdout[72] ;
wire \phy_ddio_dqdout[73] ;
wire \phy_ddio_dqdout[74] ;
wire \phy_ddio_dqdout[75] ;
wire \phy_ddio_dqdout[76] ;
wire \phy_ddio_dqdout[77] ;
wire \phy_ddio_dqdout[78] ;
wire \phy_ddio_dqdout[79] ;
wire \phy_ddio_dqdout[80] ;
wire \phy_ddio_dqdout[81] ;
wire \phy_ddio_dqdout[82] ;
wire \phy_ddio_dqdout[83] ;
wire \phy_ddio_dqdout[84] ;
wire \phy_ddio_dqdout[85] ;
wire \phy_ddio_dqdout[86] ;
wire \phy_ddio_dqdout[87] ;
wire \phy_ddio_dqdout[88] ;
wire \phy_ddio_dqdout[89] ;
wire \phy_ddio_dqdout[90] ;
wire \phy_ddio_dqdout[91] ;
wire \phy_ddio_dqdout[92] ;
wire \phy_ddio_dqdout[93] ;
wire \phy_ddio_dqdout[94] ;
wire \phy_ddio_dqdout[95] ;
wire \phy_ddio_dqdout[96] ;
wire \phy_ddio_dqdout[97] ;
wire \phy_ddio_dqdout[98] ;
wire \phy_ddio_dqdout[99] ;
wire \phy_ddio_dqdout[100] ;
wire \phy_ddio_dqdout[101] ;
wire \phy_ddio_dqdout[102] ;
wire \phy_ddio_dqdout[103] ;
wire \phy_ddio_dqdout[108] ;
wire \phy_ddio_dqdout[109] ;
wire \phy_ddio_dqdout[110] ;
wire \phy_ddio_dqdout[111] ;
wire \phy_ddio_dqdout[112] ;
wire \phy_ddio_dqdout[113] ;
wire \phy_ddio_dqdout[114] ;
wire \phy_ddio_dqdout[115] ;
wire \phy_ddio_dqdout[116] ;
wire \phy_ddio_dqdout[117] ;
wire \phy_ddio_dqdout[118] ;
wire \phy_ddio_dqdout[119] ;
wire \phy_ddio_dqdout[120] ;
wire \phy_ddio_dqdout[121] ;
wire \phy_ddio_dqdout[122] ;
wire \phy_ddio_dqdout[123] ;
wire \phy_ddio_dqdout[124] ;
wire \phy_ddio_dqdout[125] ;
wire \phy_ddio_dqdout[126] ;
wire \phy_ddio_dqdout[127] ;
wire \phy_ddio_dqdout[128] ;
wire \phy_ddio_dqdout[129] ;
wire \phy_ddio_dqdout[130] ;
wire \phy_ddio_dqdout[131] ;
wire \phy_ddio_dqdout[132] ;
wire \phy_ddio_dqdout[133] ;
wire \phy_ddio_dqdout[134] ;
wire \phy_ddio_dqdout[135] ;
wire \phy_ddio_dqdout[136] ;
wire \phy_ddio_dqdout[137] ;
wire \phy_ddio_dqdout[138] ;
wire \phy_ddio_dqdout[139] ;
wire \phy_ddio_dqoe[0] ;
wire \phy_ddio_dqoe[1] ;
wire \phy_ddio_dqoe[2] ;
wire \phy_ddio_dqoe[3] ;
wire \phy_ddio_dqoe[4] ;
wire \phy_ddio_dqoe[5] ;
wire \phy_ddio_dqoe[6] ;
wire \phy_ddio_dqoe[7] ;
wire \phy_ddio_dqoe[8] ;
wire \phy_ddio_dqoe[9] ;
wire \phy_ddio_dqoe[10] ;
wire \phy_ddio_dqoe[11] ;
wire \phy_ddio_dqoe[12] ;
wire \phy_ddio_dqoe[13] ;
wire \phy_ddio_dqoe[14] ;
wire \phy_ddio_dqoe[15] ;
wire \phy_ddio_dqoe[18] ;
wire \phy_ddio_dqoe[19] ;
wire \phy_ddio_dqoe[20] ;
wire \phy_ddio_dqoe[21] ;
wire \phy_ddio_dqoe[22] ;
wire \phy_ddio_dqoe[23] ;
wire \phy_ddio_dqoe[24] ;
wire \phy_ddio_dqoe[25] ;
wire \phy_ddio_dqoe[26] ;
wire \phy_ddio_dqoe[27] ;
wire \phy_ddio_dqoe[28] ;
wire \phy_ddio_dqoe[29] ;
wire \phy_ddio_dqoe[30] ;
wire \phy_ddio_dqoe[31] ;
wire \phy_ddio_dqoe[32] ;
wire \phy_ddio_dqoe[33] ;
wire \phy_ddio_dqoe[36] ;
wire \phy_ddio_dqoe[37] ;
wire \phy_ddio_dqoe[38] ;
wire \phy_ddio_dqoe[39] ;
wire \phy_ddio_dqoe[40] ;
wire \phy_ddio_dqoe[41] ;
wire \phy_ddio_dqoe[42] ;
wire \phy_ddio_dqoe[43] ;
wire \phy_ddio_dqoe[44] ;
wire \phy_ddio_dqoe[45] ;
wire \phy_ddio_dqoe[46] ;
wire \phy_ddio_dqoe[47] ;
wire \phy_ddio_dqoe[48] ;
wire \phy_ddio_dqoe[49] ;
wire \phy_ddio_dqoe[50] ;
wire \phy_ddio_dqoe[51] ;
wire \phy_ddio_dqoe[54] ;
wire \phy_ddio_dqoe[55] ;
wire \phy_ddio_dqoe[56] ;
wire \phy_ddio_dqoe[57] ;
wire \phy_ddio_dqoe[58] ;
wire \phy_ddio_dqoe[59] ;
wire \phy_ddio_dqoe[60] ;
wire \phy_ddio_dqoe[61] ;
wire \phy_ddio_dqoe[62] ;
wire \phy_ddio_dqoe[63] ;
wire \phy_ddio_dqoe[64] ;
wire \phy_ddio_dqoe[65] ;
wire \phy_ddio_dqoe[66] ;
wire \phy_ddio_dqoe[67] ;
wire \phy_ddio_dqoe[68] ;
wire \phy_ddio_dqoe[69] ;
wire \phy_ddio_dqs_dout[0] ;
wire \phy_ddio_dqs_dout[1] ;
wire \phy_ddio_dqs_dout[2] ;
wire \phy_ddio_dqs_dout[3] ;
wire \phy_ddio_dqs_dout[4] ;
wire \phy_ddio_dqs_dout[5] ;
wire \phy_ddio_dqs_dout[6] ;
wire \phy_ddio_dqs_dout[7] ;
wire \phy_ddio_dqs_dout[8] ;
wire \phy_ddio_dqs_dout[9] ;
wire \phy_ddio_dqs_dout[10] ;
wire \phy_ddio_dqs_dout[11] ;
wire \phy_ddio_dqs_dout[12] ;
wire \phy_ddio_dqs_dout[13] ;
wire \phy_ddio_dqs_dout[14] ;
wire \phy_ddio_dqs_dout[15] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[0] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[1] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[2] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[3] ;
wire \phy_ddio_dqslogic_aclr_pstamble[0] ;
wire \phy_ddio_dqslogic_aclr_pstamble[1] ;
wire \phy_ddio_dqslogic_aclr_pstamble[2] ;
wire \phy_ddio_dqslogic_aclr_pstamble[3] ;
wire \phy_ddio_dqslogic_dqsena[0] ;
wire \phy_ddio_dqslogic_dqsena[1] ;
wire \phy_ddio_dqslogic_dqsena[2] ;
wire \phy_ddio_dqslogic_dqsena[3] ;
wire \phy_ddio_dqslogic_dqsena[4] ;
wire \phy_ddio_dqslogic_dqsena[5] ;
wire \phy_ddio_dqslogic_dqsena[6] ;
wire \phy_ddio_dqslogic_dqsena[7] ;
wire \phy_ddio_dqslogic_fiforeset[0] ;
wire \phy_ddio_dqslogic_fiforeset[1] ;
wire \phy_ddio_dqslogic_fiforeset[2] ;
wire \phy_ddio_dqslogic_fiforeset[3] ;
wire \phy_ddio_dqslogic_incrdataen[0] ;
wire \phy_ddio_dqslogic_incrdataen[1] ;
wire \phy_ddio_dqslogic_incrdataen[2] ;
wire \phy_ddio_dqslogic_incrdataen[3] ;
wire \phy_ddio_dqslogic_incrdataen[4] ;
wire \phy_ddio_dqslogic_incrdataen[5] ;
wire \phy_ddio_dqslogic_incrdataen[6] ;
wire \phy_ddio_dqslogic_incrdataen[7] ;
wire \phy_ddio_dqslogic_incwrptr[0] ;
wire \phy_ddio_dqslogic_incwrptr[1] ;
wire \phy_ddio_dqslogic_incwrptr[2] ;
wire \phy_ddio_dqslogic_incwrptr[3] ;
wire \phy_ddio_dqslogic_incwrptr[4] ;
wire \phy_ddio_dqslogic_incwrptr[5] ;
wire \phy_ddio_dqslogic_incwrptr[6] ;
wire \phy_ddio_dqslogic_incwrptr[7] ;
wire \phy_ddio_dqslogic_oct[0] ;
wire \phy_ddio_dqslogic_oct[1] ;
wire \phy_ddio_dqslogic_oct[2] ;
wire \phy_ddio_dqslogic_oct[3] ;
wire \phy_ddio_dqslogic_oct[4] ;
wire \phy_ddio_dqslogic_oct[5] ;
wire \phy_ddio_dqslogic_oct[6] ;
wire \phy_ddio_dqslogic_oct[7] ;
wire \phy_ddio_dqslogic_readlatency[0] ;
wire \phy_ddio_dqslogic_readlatency[1] ;
wire \phy_ddio_dqslogic_readlatency[2] ;
wire \phy_ddio_dqslogic_readlatency[3] ;
wire \phy_ddio_dqslogic_readlatency[4] ;
wire \phy_ddio_dqslogic_readlatency[5] ;
wire \phy_ddio_dqslogic_readlatency[6] ;
wire \phy_ddio_dqslogic_readlatency[7] ;
wire \phy_ddio_dqslogic_readlatency[8] ;
wire \phy_ddio_dqslogic_readlatency[9] ;
wire \phy_ddio_dqslogic_readlatency[10] ;
wire \phy_ddio_dqslogic_readlatency[11] ;
wire \phy_ddio_dqslogic_readlatency[12] ;
wire \phy_ddio_dqslogic_readlatency[13] ;
wire \phy_ddio_dqslogic_readlatency[14] ;
wire \phy_ddio_dqslogic_readlatency[15] ;
wire \phy_ddio_dqslogic_readlatency[16] ;
wire \phy_ddio_dqslogic_readlatency[17] ;
wire \phy_ddio_dqslogic_readlatency[18] ;
wire \phy_ddio_dqslogic_readlatency[19] ;
wire \phy_ddio_dqs_oe[0] ;
wire \phy_ddio_dqs_oe[1] ;
wire \phy_ddio_dqs_oe[2] ;
wire \phy_ddio_dqs_oe[3] ;
wire \phy_ddio_dqs_oe[4] ;
wire \phy_ddio_dqs_oe[5] ;
wire \phy_ddio_dqs_oe[6] ;
wire \phy_ddio_dqs_oe[7] ;
wire \phy_ddio_odt[0] ;
wire \phy_ddio_odt[1] ;
wire \phy_ddio_odt[2] ;
wire \phy_ddio_odt[3] ;
wire \phy_ddio_ras_n[0] ;
wire \phy_ddio_ras_n[1] ;
wire \phy_ddio_ras_n[2] ;
wire \phy_ddio_ras_n[3] ;
wire \phy_ddio_reset_n[0] ;
wire \phy_ddio_reset_n[1] ;
wire \phy_ddio_reset_n[2] ;
wire \phy_ddio_reset_n[3] ;
wire \phy_ddio_we_n[0] ;
wire \phy_ddio_we_n[1] ;
wire \phy_ddio_we_n[2] ;
wire \phy_ddio_we_n[3] ;

wire [79:0] hphy_inst_AFIRDATA_bus;
wire [3:0] hphy_inst_AFIWLAT_bus;
wire [63:0] hphy_inst_PHYDDIOADDRDOUT_bus;
wire [11:0] hphy_inst_PHYDDIOBADOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCKDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCKEDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCSNDOUT_bus;
wire [19:0] hphy_inst_PHYDDIODMDOUT_bus;
wire [179:0] hphy_inst_PHYDDIODQDOUT_bus;
wire [89:0] hphy_inst_PHYDDIODQOE_bus;
wire [19:0] hphy_inst_PHYDDIODQSDOUT_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICDQSENA_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICFIFORESET_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICOCT_bus;
wire [24:0] hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus;
wire [9:0] hphy_inst_PHYDDIODQSOE_bus;
wire [7:0] hphy_inst_PHYDDIOODTDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORESETNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOWENDOUT_bus;

assign afi_rdata[0] = hphy_inst_AFIRDATA_bus[0];
assign afi_rdata[1] = hphy_inst_AFIRDATA_bus[1];
assign afi_rdata[2] = hphy_inst_AFIRDATA_bus[2];
assign afi_rdata[3] = hphy_inst_AFIRDATA_bus[3];
assign afi_rdata[4] = hphy_inst_AFIRDATA_bus[4];
assign afi_rdata[5] = hphy_inst_AFIRDATA_bus[5];
assign afi_rdata[6] = hphy_inst_AFIRDATA_bus[6];
assign afi_rdata[7] = hphy_inst_AFIRDATA_bus[7];
assign afi_rdata[8] = hphy_inst_AFIRDATA_bus[8];
assign afi_rdata[9] = hphy_inst_AFIRDATA_bus[9];
assign afi_rdata[10] = hphy_inst_AFIRDATA_bus[10];
assign afi_rdata[11] = hphy_inst_AFIRDATA_bus[11];
assign afi_rdata[12] = hphy_inst_AFIRDATA_bus[12];
assign afi_rdata[13] = hphy_inst_AFIRDATA_bus[13];
assign afi_rdata[14] = hphy_inst_AFIRDATA_bus[14];
assign afi_rdata[15] = hphy_inst_AFIRDATA_bus[15];
assign afi_rdata[16] = hphy_inst_AFIRDATA_bus[16];
assign afi_rdata[17] = hphy_inst_AFIRDATA_bus[17];
assign afi_rdata[18] = hphy_inst_AFIRDATA_bus[18];
assign afi_rdata[19] = hphy_inst_AFIRDATA_bus[19];
assign afi_rdata[20] = hphy_inst_AFIRDATA_bus[20];
assign afi_rdata[21] = hphy_inst_AFIRDATA_bus[21];
assign afi_rdata[22] = hphy_inst_AFIRDATA_bus[22];
assign afi_rdata[23] = hphy_inst_AFIRDATA_bus[23];
assign afi_rdata[24] = hphy_inst_AFIRDATA_bus[24];
assign afi_rdata[25] = hphy_inst_AFIRDATA_bus[25];
assign afi_rdata[26] = hphy_inst_AFIRDATA_bus[26];
assign afi_rdata[27] = hphy_inst_AFIRDATA_bus[27];
assign afi_rdata[28] = hphy_inst_AFIRDATA_bus[28];
assign afi_rdata[29] = hphy_inst_AFIRDATA_bus[29];
assign afi_rdata[30] = hphy_inst_AFIRDATA_bus[30];
assign afi_rdata[31] = hphy_inst_AFIRDATA_bus[31];
assign afi_rdata[32] = hphy_inst_AFIRDATA_bus[32];
assign afi_rdata[33] = hphy_inst_AFIRDATA_bus[33];
assign afi_rdata[34] = hphy_inst_AFIRDATA_bus[34];
assign afi_rdata[35] = hphy_inst_AFIRDATA_bus[35];
assign afi_rdata[36] = hphy_inst_AFIRDATA_bus[36];
assign afi_rdata[37] = hphy_inst_AFIRDATA_bus[37];
assign afi_rdata[38] = hphy_inst_AFIRDATA_bus[38];
assign afi_rdata[39] = hphy_inst_AFIRDATA_bus[39];
assign afi_rdata[40] = hphy_inst_AFIRDATA_bus[40];
assign afi_rdata[41] = hphy_inst_AFIRDATA_bus[41];
assign afi_rdata[42] = hphy_inst_AFIRDATA_bus[42];
assign afi_rdata[43] = hphy_inst_AFIRDATA_bus[43];
assign afi_rdata[44] = hphy_inst_AFIRDATA_bus[44];
assign afi_rdata[45] = hphy_inst_AFIRDATA_bus[45];
assign afi_rdata[46] = hphy_inst_AFIRDATA_bus[46];
assign afi_rdata[47] = hphy_inst_AFIRDATA_bus[47];
assign afi_rdata[48] = hphy_inst_AFIRDATA_bus[48];
assign afi_rdata[49] = hphy_inst_AFIRDATA_bus[49];
assign afi_rdata[50] = hphy_inst_AFIRDATA_bus[50];
assign afi_rdata[51] = hphy_inst_AFIRDATA_bus[51];
assign afi_rdata[52] = hphy_inst_AFIRDATA_bus[52];
assign afi_rdata[53] = hphy_inst_AFIRDATA_bus[53];
assign afi_rdata[54] = hphy_inst_AFIRDATA_bus[54];
assign afi_rdata[55] = hphy_inst_AFIRDATA_bus[55];
assign afi_rdata[56] = hphy_inst_AFIRDATA_bus[56];
assign afi_rdata[57] = hphy_inst_AFIRDATA_bus[57];
assign afi_rdata[58] = hphy_inst_AFIRDATA_bus[58];
assign afi_rdata[59] = hphy_inst_AFIRDATA_bus[59];
assign afi_rdata[60] = hphy_inst_AFIRDATA_bus[60];
assign afi_rdata[61] = hphy_inst_AFIRDATA_bus[61];
assign afi_rdata[62] = hphy_inst_AFIRDATA_bus[62];
assign afi_rdata[63] = hphy_inst_AFIRDATA_bus[63];
assign afi_rdata[64] = hphy_inst_AFIRDATA_bus[64];
assign afi_rdata[65] = hphy_inst_AFIRDATA_bus[65];
assign afi_rdata[66] = hphy_inst_AFIRDATA_bus[66];
assign afi_rdata[67] = hphy_inst_AFIRDATA_bus[67];
assign afi_rdata[68] = hphy_inst_AFIRDATA_bus[68];
assign afi_rdata[69] = hphy_inst_AFIRDATA_bus[69];
assign afi_rdata[70] = hphy_inst_AFIRDATA_bus[70];
assign afi_rdata[71] = hphy_inst_AFIRDATA_bus[71];
assign afi_rdata[72] = hphy_inst_AFIRDATA_bus[72];
assign afi_rdata[73] = hphy_inst_AFIRDATA_bus[73];
assign afi_rdata[74] = hphy_inst_AFIRDATA_bus[74];
assign afi_rdata[75] = hphy_inst_AFIRDATA_bus[75];
assign afi_rdata[76] = hphy_inst_AFIRDATA_bus[76];
assign afi_rdata[77] = hphy_inst_AFIRDATA_bus[77];
assign afi_rdata[78] = hphy_inst_AFIRDATA_bus[78];
assign afi_rdata[79] = hphy_inst_AFIRDATA_bus[79];

assign afi_wlat[0] = hphy_inst_AFIWLAT_bus[0];
assign afi_wlat[1] = hphy_inst_AFIWLAT_bus[1];
assign afi_wlat[2] = hphy_inst_AFIWLAT_bus[2];
assign afi_wlat[3] = hphy_inst_AFIWLAT_bus[3];

assign \phy_ddio_address[0]  = hphy_inst_PHYDDIOADDRDOUT_bus[0];
assign \phy_ddio_address[1]  = hphy_inst_PHYDDIOADDRDOUT_bus[1];
assign \phy_ddio_address[2]  = hphy_inst_PHYDDIOADDRDOUT_bus[2];
assign \phy_ddio_address[3]  = hphy_inst_PHYDDIOADDRDOUT_bus[3];
assign \phy_ddio_address[4]  = hphy_inst_PHYDDIOADDRDOUT_bus[4];
assign \phy_ddio_address[5]  = hphy_inst_PHYDDIOADDRDOUT_bus[5];
assign \phy_ddio_address[6]  = hphy_inst_PHYDDIOADDRDOUT_bus[6];
assign \phy_ddio_address[7]  = hphy_inst_PHYDDIOADDRDOUT_bus[7];
assign \phy_ddio_address[8]  = hphy_inst_PHYDDIOADDRDOUT_bus[8];
assign \phy_ddio_address[9]  = hphy_inst_PHYDDIOADDRDOUT_bus[9];
assign \phy_ddio_address[10]  = hphy_inst_PHYDDIOADDRDOUT_bus[10];
assign \phy_ddio_address[11]  = hphy_inst_PHYDDIOADDRDOUT_bus[11];
assign \phy_ddio_address[12]  = hphy_inst_PHYDDIOADDRDOUT_bus[12];
assign \phy_ddio_address[13]  = hphy_inst_PHYDDIOADDRDOUT_bus[13];
assign \phy_ddio_address[14]  = hphy_inst_PHYDDIOADDRDOUT_bus[14];
assign \phy_ddio_address[15]  = hphy_inst_PHYDDIOADDRDOUT_bus[15];
assign \phy_ddio_address[16]  = hphy_inst_PHYDDIOADDRDOUT_bus[16];
assign \phy_ddio_address[17]  = hphy_inst_PHYDDIOADDRDOUT_bus[17];
assign \phy_ddio_address[18]  = hphy_inst_PHYDDIOADDRDOUT_bus[18];
assign \phy_ddio_address[19]  = hphy_inst_PHYDDIOADDRDOUT_bus[19];
assign \phy_ddio_address[20]  = hphy_inst_PHYDDIOADDRDOUT_bus[20];
assign \phy_ddio_address[21]  = hphy_inst_PHYDDIOADDRDOUT_bus[21];
assign \phy_ddio_address[22]  = hphy_inst_PHYDDIOADDRDOUT_bus[22];
assign \phy_ddio_address[23]  = hphy_inst_PHYDDIOADDRDOUT_bus[23];
assign \phy_ddio_address[24]  = hphy_inst_PHYDDIOADDRDOUT_bus[24];
assign \phy_ddio_address[25]  = hphy_inst_PHYDDIOADDRDOUT_bus[25];
assign \phy_ddio_address[26]  = hphy_inst_PHYDDIOADDRDOUT_bus[26];
assign \phy_ddio_address[27]  = hphy_inst_PHYDDIOADDRDOUT_bus[27];
assign \phy_ddio_address[28]  = hphy_inst_PHYDDIOADDRDOUT_bus[28];
assign \phy_ddio_address[29]  = hphy_inst_PHYDDIOADDRDOUT_bus[29];
assign \phy_ddio_address[30]  = hphy_inst_PHYDDIOADDRDOUT_bus[30];
assign \phy_ddio_address[31]  = hphy_inst_PHYDDIOADDRDOUT_bus[31];
assign \phy_ddio_address[32]  = hphy_inst_PHYDDIOADDRDOUT_bus[32];
assign \phy_ddio_address[33]  = hphy_inst_PHYDDIOADDRDOUT_bus[33];
assign \phy_ddio_address[34]  = hphy_inst_PHYDDIOADDRDOUT_bus[34];
assign \phy_ddio_address[35]  = hphy_inst_PHYDDIOADDRDOUT_bus[35];
assign \phy_ddio_address[36]  = hphy_inst_PHYDDIOADDRDOUT_bus[36];
assign \phy_ddio_address[37]  = hphy_inst_PHYDDIOADDRDOUT_bus[37];
assign \phy_ddio_address[38]  = hphy_inst_PHYDDIOADDRDOUT_bus[38];
assign \phy_ddio_address[39]  = hphy_inst_PHYDDIOADDRDOUT_bus[39];
assign \phy_ddio_address[40]  = hphy_inst_PHYDDIOADDRDOUT_bus[40];
assign \phy_ddio_address[41]  = hphy_inst_PHYDDIOADDRDOUT_bus[41];
assign \phy_ddio_address[42]  = hphy_inst_PHYDDIOADDRDOUT_bus[42];
assign \phy_ddio_address[43]  = hphy_inst_PHYDDIOADDRDOUT_bus[43];
assign \phy_ddio_address[44]  = hphy_inst_PHYDDIOADDRDOUT_bus[44];
assign \phy_ddio_address[45]  = hphy_inst_PHYDDIOADDRDOUT_bus[45];
assign \phy_ddio_address[46]  = hphy_inst_PHYDDIOADDRDOUT_bus[46];
assign \phy_ddio_address[47]  = hphy_inst_PHYDDIOADDRDOUT_bus[47];
assign \phy_ddio_address[48]  = hphy_inst_PHYDDIOADDRDOUT_bus[48];
assign \phy_ddio_address[49]  = hphy_inst_PHYDDIOADDRDOUT_bus[49];
assign \phy_ddio_address[50]  = hphy_inst_PHYDDIOADDRDOUT_bus[50];
assign \phy_ddio_address[51]  = hphy_inst_PHYDDIOADDRDOUT_bus[51];
assign \phy_ddio_address[52]  = hphy_inst_PHYDDIOADDRDOUT_bus[52];
assign \phy_ddio_address[53]  = hphy_inst_PHYDDIOADDRDOUT_bus[53];
assign \phy_ddio_address[54]  = hphy_inst_PHYDDIOADDRDOUT_bus[54];
assign \phy_ddio_address[55]  = hphy_inst_PHYDDIOADDRDOUT_bus[55];
assign \phy_ddio_address[56]  = hphy_inst_PHYDDIOADDRDOUT_bus[56];
assign \phy_ddio_address[57]  = hphy_inst_PHYDDIOADDRDOUT_bus[57];
assign \phy_ddio_address[58]  = hphy_inst_PHYDDIOADDRDOUT_bus[58];
assign \phy_ddio_address[59]  = hphy_inst_PHYDDIOADDRDOUT_bus[59];

assign \phy_ddio_bank[0]  = hphy_inst_PHYDDIOBADOUT_bus[0];
assign \phy_ddio_bank[1]  = hphy_inst_PHYDDIOBADOUT_bus[1];
assign \phy_ddio_bank[2]  = hphy_inst_PHYDDIOBADOUT_bus[2];
assign \phy_ddio_bank[3]  = hphy_inst_PHYDDIOBADOUT_bus[3];
assign \phy_ddio_bank[4]  = hphy_inst_PHYDDIOBADOUT_bus[4];
assign \phy_ddio_bank[5]  = hphy_inst_PHYDDIOBADOUT_bus[5];
assign \phy_ddio_bank[6]  = hphy_inst_PHYDDIOBADOUT_bus[6];
assign \phy_ddio_bank[7]  = hphy_inst_PHYDDIOBADOUT_bus[7];
assign \phy_ddio_bank[8]  = hphy_inst_PHYDDIOBADOUT_bus[8];
assign \phy_ddio_bank[9]  = hphy_inst_PHYDDIOBADOUT_bus[9];
assign \phy_ddio_bank[10]  = hphy_inst_PHYDDIOBADOUT_bus[10];
assign \phy_ddio_bank[11]  = hphy_inst_PHYDDIOBADOUT_bus[11];

assign \phy_ddio_cas_n[0]  = hphy_inst_PHYDDIOCASNDOUT_bus[0];
assign \phy_ddio_cas_n[1]  = hphy_inst_PHYDDIOCASNDOUT_bus[1];
assign \phy_ddio_cas_n[2]  = hphy_inst_PHYDDIOCASNDOUT_bus[2];
assign \phy_ddio_cas_n[3]  = hphy_inst_PHYDDIOCASNDOUT_bus[3];

assign \phy_ddio_ck[0]  = hphy_inst_PHYDDIOCKDOUT_bus[0];
assign \phy_ddio_ck[1]  = hphy_inst_PHYDDIOCKDOUT_bus[1];

assign \phy_ddio_cke[0]  = hphy_inst_PHYDDIOCKEDOUT_bus[0];
assign \phy_ddio_cke[1]  = hphy_inst_PHYDDIOCKEDOUT_bus[1];
assign \phy_ddio_cke[2]  = hphy_inst_PHYDDIOCKEDOUT_bus[2];
assign \phy_ddio_cke[3]  = hphy_inst_PHYDDIOCKEDOUT_bus[3];

assign \phy_ddio_cs_n[0]  = hphy_inst_PHYDDIOCSNDOUT_bus[0];
assign \phy_ddio_cs_n[1]  = hphy_inst_PHYDDIOCSNDOUT_bus[1];
assign \phy_ddio_cs_n[2]  = hphy_inst_PHYDDIOCSNDOUT_bus[2];
assign \phy_ddio_cs_n[3]  = hphy_inst_PHYDDIOCSNDOUT_bus[3];

assign \phy_ddio_dmdout[0]  = hphy_inst_PHYDDIODMDOUT_bus[0];
assign \phy_ddio_dmdout[1]  = hphy_inst_PHYDDIODMDOUT_bus[1];
assign \phy_ddio_dmdout[2]  = hphy_inst_PHYDDIODMDOUT_bus[2];
assign \phy_ddio_dmdout[3]  = hphy_inst_PHYDDIODMDOUT_bus[3];
assign \phy_ddio_dmdout[4]  = hphy_inst_PHYDDIODMDOUT_bus[4];
assign \phy_ddio_dmdout[5]  = hphy_inst_PHYDDIODMDOUT_bus[5];
assign \phy_ddio_dmdout[6]  = hphy_inst_PHYDDIODMDOUT_bus[6];
assign \phy_ddio_dmdout[7]  = hphy_inst_PHYDDIODMDOUT_bus[7];
assign \phy_ddio_dmdout[8]  = hphy_inst_PHYDDIODMDOUT_bus[8];
assign \phy_ddio_dmdout[9]  = hphy_inst_PHYDDIODMDOUT_bus[9];
assign \phy_ddio_dmdout[10]  = hphy_inst_PHYDDIODMDOUT_bus[10];
assign \phy_ddio_dmdout[11]  = hphy_inst_PHYDDIODMDOUT_bus[11];
assign \phy_ddio_dmdout[12]  = hphy_inst_PHYDDIODMDOUT_bus[12];
assign \phy_ddio_dmdout[13]  = hphy_inst_PHYDDIODMDOUT_bus[13];
assign \phy_ddio_dmdout[14]  = hphy_inst_PHYDDIODMDOUT_bus[14];
assign \phy_ddio_dmdout[15]  = hphy_inst_PHYDDIODMDOUT_bus[15];

assign \phy_ddio_dqdout[0]  = hphy_inst_PHYDDIODQDOUT_bus[0];
assign \phy_ddio_dqdout[1]  = hphy_inst_PHYDDIODQDOUT_bus[1];
assign \phy_ddio_dqdout[2]  = hphy_inst_PHYDDIODQDOUT_bus[2];
assign \phy_ddio_dqdout[3]  = hphy_inst_PHYDDIODQDOUT_bus[3];
assign \phy_ddio_dqdout[4]  = hphy_inst_PHYDDIODQDOUT_bus[4];
assign \phy_ddio_dqdout[5]  = hphy_inst_PHYDDIODQDOUT_bus[5];
assign \phy_ddio_dqdout[6]  = hphy_inst_PHYDDIODQDOUT_bus[6];
assign \phy_ddio_dqdout[7]  = hphy_inst_PHYDDIODQDOUT_bus[7];
assign \phy_ddio_dqdout[8]  = hphy_inst_PHYDDIODQDOUT_bus[8];
assign \phy_ddio_dqdout[9]  = hphy_inst_PHYDDIODQDOUT_bus[9];
assign \phy_ddio_dqdout[10]  = hphy_inst_PHYDDIODQDOUT_bus[10];
assign \phy_ddio_dqdout[11]  = hphy_inst_PHYDDIODQDOUT_bus[11];
assign \phy_ddio_dqdout[12]  = hphy_inst_PHYDDIODQDOUT_bus[12];
assign \phy_ddio_dqdout[13]  = hphy_inst_PHYDDIODQDOUT_bus[13];
assign \phy_ddio_dqdout[14]  = hphy_inst_PHYDDIODQDOUT_bus[14];
assign \phy_ddio_dqdout[15]  = hphy_inst_PHYDDIODQDOUT_bus[15];
assign \phy_ddio_dqdout[16]  = hphy_inst_PHYDDIODQDOUT_bus[16];
assign \phy_ddio_dqdout[17]  = hphy_inst_PHYDDIODQDOUT_bus[17];
assign \phy_ddio_dqdout[18]  = hphy_inst_PHYDDIODQDOUT_bus[18];
assign \phy_ddio_dqdout[19]  = hphy_inst_PHYDDIODQDOUT_bus[19];
assign \phy_ddio_dqdout[20]  = hphy_inst_PHYDDIODQDOUT_bus[20];
assign \phy_ddio_dqdout[21]  = hphy_inst_PHYDDIODQDOUT_bus[21];
assign \phy_ddio_dqdout[22]  = hphy_inst_PHYDDIODQDOUT_bus[22];
assign \phy_ddio_dqdout[23]  = hphy_inst_PHYDDIODQDOUT_bus[23];
assign \phy_ddio_dqdout[24]  = hphy_inst_PHYDDIODQDOUT_bus[24];
assign \phy_ddio_dqdout[25]  = hphy_inst_PHYDDIODQDOUT_bus[25];
assign \phy_ddio_dqdout[26]  = hphy_inst_PHYDDIODQDOUT_bus[26];
assign \phy_ddio_dqdout[27]  = hphy_inst_PHYDDIODQDOUT_bus[27];
assign \phy_ddio_dqdout[28]  = hphy_inst_PHYDDIODQDOUT_bus[28];
assign \phy_ddio_dqdout[29]  = hphy_inst_PHYDDIODQDOUT_bus[29];
assign \phy_ddio_dqdout[30]  = hphy_inst_PHYDDIODQDOUT_bus[30];
assign \phy_ddio_dqdout[31]  = hphy_inst_PHYDDIODQDOUT_bus[31];
assign \phy_ddio_dqdout[36]  = hphy_inst_PHYDDIODQDOUT_bus[36];
assign \phy_ddio_dqdout[37]  = hphy_inst_PHYDDIODQDOUT_bus[37];
assign \phy_ddio_dqdout[38]  = hphy_inst_PHYDDIODQDOUT_bus[38];
assign \phy_ddio_dqdout[39]  = hphy_inst_PHYDDIODQDOUT_bus[39];
assign \phy_ddio_dqdout[40]  = hphy_inst_PHYDDIODQDOUT_bus[40];
assign \phy_ddio_dqdout[41]  = hphy_inst_PHYDDIODQDOUT_bus[41];
assign \phy_ddio_dqdout[42]  = hphy_inst_PHYDDIODQDOUT_bus[42];
assign \phy_ddio_dqdout[43]  = hphy_inst_PHYDDIODQDOUT_bus[43];
assign \phy_ddio_dqdout[44]  = hphy_inst_PHYDDIODQDOUT_bus[44];
assign \phy_ddio_dqdout[45]  = hphy_inst_PHYDDIODQDOUT_bus[45];
assign \phy_ddio_dqdout[46]  = hphy_inst_PHYDDIODQDOUT_bus[46];
assign \phy_ddio_dqdout[47]  = hphy_inst_PHYDDIODQDOUT_bus[47];
assign \phy_ddio_dqdout[48]  = hphy_inst_PHYDDIODQDOUT_bus[48];
assign \phy_ddio_dqdout[49]  = hphy_inst_PHYDDIODQDOUT_bus[49];
assign \phy_ddio_dqdout[50]  = hphy_inst_PHYDDIODQDOUT_bus[50];
assign \phy_ddio_dqdout[51]  = hphy_inst_PHYDDIODQDOUT_bus[51];
assign \phy_ddio_dqdout[52]  = hphy_inst_PHYDDIODQDOUT_bus[52];
assign \phy_ddio_dqdout[53]  = hphy_inst_PHYDDIODQDOUT_bus[53];
assign \phy_ddio_dqdout[54]  = hphy_inst_PHYDDIODQDOUT_bus[54];
assign \phy_ddio_dqdout[55]  = hphy_inst_PHYDDIODQDOUT_bus[55];
assign \phy_ddio_dqdout[56]  = hphy_inst_PHYDDIODQDOUT_bus[56];
assign \phy_ddio_dqdout[57]  = hphy_inst_PHYDDIODQDOUT_bus[57];
assign \phy_ddio_dqdout[58]  = hphy_inst_PHYDDIODQDOUT_bus[58];
assign \phy_ddio_dqdout[59]  = hphy_inst_PHYDDIODQDOUT_bus[59];
assign \phy_ddio_dqdout[60]  = hphy_inst_PHYDDIODQDOUT_bus[60];
assign \phy_ddio_dqdout[61]  = hphy_inst_PHYDDIODQDOUT_bus[61];
assign \phy_ddio_dqdout[62]  = hphy_inst_PHYDDIODQDOUT_bus[62];
assign \phy_ddio_dqdout[63]  = hphy_inst_PHYDDIODQDOUT_bus[63];
assign \phy_ddio_dqdout[64]  = hphy_inst_PHYDDIODQDOUT_bus[64];
assign \phy_ddio_dqdout[65]  = hphy_inst_PHYDDIODQDOUT_bus[65];
assign \phy_ddio_dqdout[66]  = hphy_inst_PHYDDIODQDOUT_bus[66];
assign \phy_ddio_dqdout[67]  = hphy_inst_PHYDDIODQDOUT_bus[67];
assign \phy_ddio_dqdout[72]  = hphy_inst_PHYDDIODQDOUT_bus[72];
assign \phy_ddio_dqdout[73]  = hphy_inst_PHYDDIODQDOUT_bus[73];
assign \phy_ddio_dqdout[74]  = hphy_inst_PHYDDIODQDOUT_bus[74];
assign \phy_ddio_dqdout[75]  = hphy_inst_PHYDDIODQDOUT_bus[75];
assign \phy_ddio_dqdout[76]  = hphy_inst_PHYDDIODQDOUT_bus[76];
assign \phy_ddio_dqdout[77]  = hphy_inst_PHYDDIODQDOUT_bus[77];
assign \phy_ddio_dqdout[78]  = hphy_inst_PHYDDIODQDOUT_bus[78];
assign \phy_ddio_dqdout[79]  = hphy_inst_PHYDDIODQDOUT_bus[79];
assign \phy_ddio_dqdout[80]  = hphy_inst_PHYDDIODQDOUT_bus[80];
assign \phy_ddio_dqdout[81]  = hphy_inst_PHYDDIODQDOUT_bus[81];
assign \phy_ddio_dqdout[82]  = hphy_inst_PHYDDIODQDOUT_bus[82];
assign \phy_ddio_dqdout[83]  = hphy_inst_PHYDDIODQDOUT_bus[83];
assign \phy_ddio_dqdout[84]  = hphy_inst_PHYDDIODQDOUT_bus[84];
assign \phy_ddio_dqdout[85]  = hphy_inst_PHYDDIODQDOUT_bus[85];
assign \phy_ddio_dqdout[86]  = hphy_inst_PHYDDIODQDOUT_bus[86];
assign \phy_ddio_dqdout[87]  = hphy_inst_PHYDDIODQDOUT_bus[87];
assign \phy_ddio_dqdout[88]  = hphy_inst_PHYDDIODQDOUT_bus[88];
assign \phy_ddio_dqdout[89]  = hphy_inst_PHYDDIODQDOUT_bus[89];
assign \phy_ddio_dqdout[90]  = hphy_inst_PHYDDIODQDOUT_bus[90];
assign \phy_ddio_dqdout[91]  = hphy_inst_PHYDDIODQDOUT_bus[91];
assign \phy_ddio_dqdout[92]  = hphy_inst_PHYDDIODQDOUT_bus[92];
assign \phy_ddio_dqdout[93]  = hphy_inst_PHYDDIODQDOUT_bus[93];
assign \phy_ddio_dqdout[94]  = hphy_inst_PHYDDIODQDOUT_bus[94];
assign \phy_ddio_dqdout[95]  = hphy_inst_PHYDDIODQDOUT_bus[95];
assign \phy_ddio_dqdout[96]  = hphy_inst_PHYDDIODQDOUT_bus[96];
assign \phy_ddio_dqdout[97]  = hphy_inst_PHYDDIODQDOUT_bus[97];
assign \phy_ddio_dqdout[98]  = hphy_inst_PHYDDIODQDOUT_bus[98];
assign \phy_ddio_dqdout[99]  = hphy_inst_PHYDDIODQDOUT_bus[99];
assign \phy_ddio_dqdout[100]  = hphy_inst_PHYDDIODQDOUT_bus[100];
assign \phy_ddio_dqdout[101]  = hphy_inst_PHYDDIODQDOUT_bus[101];
assign \phy_ddio_dqdout[102]  = hphy_inst_PHYDDIODQDOUT_bus[102];
assign \phy_ddio_dqdout[103]  = hphy_inst_PHYDDIODQDOUT_bus[103];
assign \phy_ddio_dqdout[108]  = hphy_inst_PHYDDIODQDOUT_bus[108];
assign \phy_ddio_dqdout[109]  = hphy_inst_PHYDDIODQDOUT_bus[109];
assign \phy_ddio_dqdout[110]  = hphy_inst_PHYDDIODQDOUT_bus[110];
assign \phy_ddio_dqdout[111]  = hphy_inst_PHYDDIODQDOUT_bus[111];
assign \phy_ddio_dqdout[112]  = hphy_inst_PHYDDIODQDOUT_bus[112];
assign \phy_ddio_dqdout[113]  = hphy_inst_PHYDDIODQDOUT_bus[113];
assign \phy_ddio_dqdout[114]  = hphy_inst_PHYDDIODQDOUT_bus[114];
assign \phy_ddio_dqdout[115]  = hphy_inst_PHYDDIODQDOUT_bus[115];
assign \phy_ddio_dqdout[116]  = hphy_inst_PHYDDIODQDOUT_bus[116];
assign \phy_ddio_dqdout[117]  = hphy_inst_PHYDDIODQDOUT_bus[117];
assign \phy_ddio_dqdout[118]  = hphy_inst_PHYDDIODQDOUT_bus[118];
assign \phy_ddio_dqdout[119]  = hphy_inst_PHYDDIODQDOUT_bus[119];
assign \phy_ddio_dqdout[120]  = hphy_inst_PHYDDIODQDOUT_bus[120];
assign \phy_ddio_dqdout[121]  = hphy_inst_PHYDDIODQDOUT_bus[121];
assign \phy_ddio_dqdout[122]  = hphy_inst_PHYDDIODQDOUT_bus[122];
assign \phy_ddio_dqdout[123]  = hphy_inst_PHYDDIODQDOUT_bus[123];
assign \phy_ddio_dqdout[124]  = hphy_inst_PHYDDIODQDOUT_bus[124];
assign \phy_ddio_dqdout[125]  = hphy_inst_PHYDDIODQDOUT_bus[125];
assign \phy_ddio_dqdout[126]  = hphy_inst_PHYDDIODQDOUT_bus[126];
assign \phy_ddio_dqdout[127]  = hphy_inst_PHYDDIODQDOUT_bus[127];
assign \phy_ddio_dqdout[128]  = hphy_inst_PHYDDIODQDOUT_bus[128];
assign \phy_ddio_dqdout[129]  = hphy_inst_PHYDDIODQDOUT_bus[129];
assign \phy_ddio_dqdout[130]  = hphy_inst_PHYDDIODQDOUT_bus[130];
assign \phy_ddio_dqdout[131]  = hphy_inst_PHYDDIODQDOUT_bus[131];
assign \phy_ddio_dqdout[132]  = hphy_inst_PHYDDIODQDOUT_bus[132];
assign \phy_ddio_dqdout[133]  = hphy_inst_PHYDDIODQDOUT_bus[133];
assign \phy_ddio_dqdout[134]  = hphy_inst_PHYDDIODQDOUT_bus[134];
assign \phy_ddio_dqdout[135]  = hphy_inst_PHYDDIODQDOUT_bus[135];
assign \phy_ddio_dqdout[136]  = hphy_inst_PHYDDIODQDOUT_bus[136];
assign \phy_ddio_dqdout[137]  = hphy_inst_PHYDDIODQDOUT_bus[137];
assign \phy_ddio_dqdout[138]  = hphy_inst_PHYDDIODQDOUT_bus[138];
assign \phy_ddio_dqdout[139]  = hphy_inst_PHYDDIODQDOUT_bus[139];

assign \phy_ddio_dqoe[0]  = hphy_inst_PHYDDIODQOE_bus[0];
assign \phy_ddio_dqoe[1]  = hphy_inst_PHYDDIODQOE_bus[1];
assign \phy_ddio_dqoe[2]  = hphy_inst_PHYDDIODQOE_bus[2];
assign \phy_ddio_dqoe[3]  = hphy_inst_PHYDDIODQOE_bus[3];
assign \phy_ddio_dqoe[4]  = hphy_inst_PHYDDIODQOE_bus[4];
assign \phy_ddio_dqoe[5]  = hphy_inst_PHYDDIODQOE_bus[5];
assign \phy_ddio_dqoe[6]  = hphy_inst_PHYDDIODQOE_bus[6];
assign \phy_ddio_dqoe[7]  = hphy_inst_PHYDDIODQOE_bus[7];
assign \phy_ddio_dqoe[8]  = hphy_inst_PHYDDIODQOE_bus[8];
assign \phy_ddio_dqoe[9]  = hphy_inst_PHYDDIODQOE_bus[9];
assign \phy_ddio_dqoe[10]  = hphy_inst_PHYDDIODQOE_bus[10];
assign \phy_ddio_dqoe[11]  = hphy_inst_PHYDDIODQOE_bus[11];
assign \phy_ddio_dqoe[12]  = hphy_inst_PHYDDIODQOE_bus[12];
assign \phy_ddio_dqoe[13]  = hphy_inst_PHYDDIODQOE_bus[13];
assign \phy_ddio_dqoe[14]  = hphy_inst_PHYDDIODQOE_bus[14];
assign \phy_ddio_dqoe[15]  = hphy_inst_PHYDDIODQOE_bus[15];
assign \phy_ddio_dqoe[18]  = hphy_inst_PHYDDIODQOE_bus[18];
assign \phy_ddio_dqoe[19]  = hphy_inst_PHYDDIODQOE_bus[19];
assign \phy_ddio_dqoe[20]  = hphy_inst_PHYDDIODQOE_bus[20];
assign \phy_ddio_dqoe[21]  = hphy_inst_PHYDDIODQOE_bus[21];
assign \phy_ddio_dqoe[22]  = hphy_inst_PHYDDIODQOE_bus[22];
assign \phy_ddio_dqoe[23]  = hphy_inst_PHYDDIODQOE_bus[23];
assign \phy_ddio_dqoe[24]  = hphy_inst_PHYDDIODQOE_bus[24];
assign \phy_ddio_dqoe[25]  = hphy_inst_PHYDDIODQOE_bus[25];
assign \phy_ddio_dqoe[26]  = hphy_inst_PHYDDIODQOE_bus[26];
assign \phy_ddio_dqoe[27]  = hphy_inst_PHYDDIODQOE_bus[27];
assign \phy_ddio_dqoe[28]  = hphy_inst_PHYDDIODQOE_bus[28];
assign \phy_ddio_dqoe[29]  = hphy_inst_PHYDDIODQOE_bus[29];
assign \phy_ddio_dqoe[30]  = hphy_inst_PHYDDIODQOE_bus[30];
assign \phy_ddio_dqoe[31]  = hphy_inst_PHYDDIODQOE_bus[31];
assign \phy_ddio_dqoe[32]  = hphy_inst_PHYDDIODQOE_bus[32];
assign \phy_ddio_dqoe[33]  = hphy_inst_PHYDDIODQOE_bus[33];
assign \phy_ddio_dqoe[36]  = hphy_inst_PHYDDIODQOE_bus[36];
assign \phy_ddio_dqoe[37]  = hphy_inst_PHYDDIODQOE_bus[37];
assign \phy_ddio_dqoe[38]  = hphy_inst_PHYDDIODQOE_bus[38];
assign \phy_ddio_dqoe[39]  = hphy_inst_PHYDDIODQOE_bus[39];
assign \phy_ddio_dqoe[40]  = hphy_inst_PHYDDIODQOE_bus[40];
assign \phy_ddio_dqoe[41]  = hphy_inst_PHYDDIODQOE_bus[41];
assign \phy_ddio_dqoe[42]  = hphy_inst_PHYDDIODQOE_bus[42];
assign \phy_ddio_dqoe[43]  = hphy_inst_PHYDDIODQOE_bus[43];
assign \phy_ddio_dqoe[44]  = hphy_inst_PHYDDIODQOE_bus[44];
assign \phy_ddio_dqoe[45]  = hphy_inst_PHYDDIODQOE_bus[45];
assign \phy_ddio_dqoe[46]  = hphy_inst_PHYDDIODQOE_bus[46];
assign \phy_ddio_dqoe[47]  = hphy_inst_PHYDDIODQOE_bus[47];
assign \phy_ddio_dqoe[48]  = hphy_inst_PHYDDIODQOE_bus[48];
assign \phy_ddio_dqoe[49]  = hphy_inst_PHYDDIODQOE_bus[49];
assign \phy_ddio_dqoe[50]  = hphy_inst_PHYDDIODQOE_bus[50];
assign \phy_ddio_dqoe[51]  = hphy_inst_PHYDDIODQOE_bus[51];
assign \phy_ddio_dqoe[54]  = hphy_inst_PHYDDIODQOE_bus[54];
assign \phy_ddio_dqoe[55]  = hphy_inst_PHYDDIODQOE_bus[55];
assign \phy_ddio_dqoe[56]  = hphy_inst_PHYDDIODQOE_bus[56];
assign \phy_ddio_dqoe[57]  = hphy_inst_PHYDDIODQOE_bus[57];
assign \phy_ddio_dqoe[58]  = hphy_inst_PHYDDIODQOE_bus[58];
assign \phy_ddio_dqoe[59]  = hphy_inst_PHYDDIODQOE_bus[59];
assign \phy_ddio_dqoe[60]  = hphy_inst_PHYDDIODQOE_bus[60];
assign \phy_ddio_dqoe[61]  = hphy_inst_PHYDDIODQOE_bus[61];
assign \phy_ddio_dqoe[62]  = hphy_inst_PHYDDIODQOE_bus[62];
assign \phy_ddio_dqoe[63]  = hphy_inst_PHYDDIODQOE_bus[63];
assign \phy_ddio_dqoe[64]  = hphy_inst_PHYDDIODQOE_bus[64];
assign \phy_ddio_dqoe[65]  = hphy_inst_PHYDDIODQOE_bus[65];
assign \phy_ddio_dqoe[66]  = hphy_inst_PHYDDIODQOE_bus[66];
assign \phy_ddio_dqoe[67]  = hphy_inst_PHYDDIODQOE_bus[67];
assign \phy_ddio_dqoe[68]  = hphy_inst_PHYDDIODQOE_bus[68];
assign \phy_ddio_dqoe[69]  = hphy_inst_PHYDDIODQOE_bus[69];

assign \phy_ddio_dqs_dout[0]  = hphy_inst_PHYDDIODQSDOUT_bus[0];
assign \phy_ddio_dqs_dout[1]  = hphy_inst_PHYDDIODQSDOUT_bus[1];
assign \phy_ddio_dqs_dout[2]  = hphy_inst_PHYDDIODQSDOUT_bus[2];
assign \phy_ddio_dqs_dout[3]  = hphy_inst_PHYDDIODQSDOUT_bus[3];
assign \phy_ddio_dqs_dout[4]  = hphy_inst_PHYDDIODQSDOUT_bus[4];
assign \phy_ddio_dqs_dout[5]  = hphy_inst_PHYDDIODQSDOUT_bus[5];
assign \phy_ddio_dqs_dout[6]  = hphy_inst_PHYDDIODQSDOUT_bus[6];
assign \phy_ddio_dqs_dout[7]  = hphy_inst_PHYDDIODQSDOUT_bus[7];
assign \phy_ddio_dqs_dout[8]  = hphy_inst_PHYDDIODQSDOUT_bus[8];
assign \phy_ddio_dqs_dout[9]  = hphy_inst_PHYDDIODQSDOUT_bus[9];
assign \phy_ddio_dqs_dout[10]  = hphy_inst_PHYDDIODQSDOUT_bus[10];
assign \phy_ddio_dqs_dout[11]  = hphy_inst_PHYDDIODQSDOUT_bus[11];
assign \phy_ddio_dqs_dout[12]  = hphy_inst_PHYDDIODQSDOUT_bus[12];
assign \phy_ddio_dqs_dout[13]  = hphy_inst_PHYDDIODQSDOUT_bus[13];
assign \phy_ddio_dqs_dout[14]  = hphy_inst_PHYDDIODQSDOUT_bus[14];
assign \phy_ddio_dqs_dout[15]  = hphy_inst_PHYDDIODQSDOUT_bus[15];

assign \phy_ddio_dqslogic_aclr_fifoctrl[0]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[0];
assign \phy_ddio_dqslogic_aclr_fifoctrl[1]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[1];
assign \phy_ddio_dqslogic_aclr_fifoctrl[2]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[2];
assign \phy_ddio_dqslogic_aclr_fifoctrl[3]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[3];

assign \phy_ddio_dqslogic_aclr_pstamble[0]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[0];
assign \phy_ddio_dqslogic_aclr_pstamble[1]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[1];
assign \phy_ddio_dqslogic_aclr_pstamble[2]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[2];
assign \phy_ddio_dqslogic_aclr_pstamble[3]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[3];

assign \phy_ddio_dqslogic_dqsena[0]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[0];
assign \phy_ddio_dqslogic_dqsena[1]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[1];
assign \phy_ddio_dqslogic_dqsena[2]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[2];
assign \phy_ddio_dqslogic_dqsena[3]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[3];
assign \phy_ddio_dqslogic_dqsena[4]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[4];
assign \phy_ddio_dqslogic_dqsena[5]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[5];
assign \phy_ddio_dqslogic_dqsena[6]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[6];
assign \phy_ddio_dqslogic_dqsena[7]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[7];

assign \phy_ddio_dqslogic_fiforeset[0]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[0];
assign \phy_ddio_dqslogic_fiforeset[1]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[1];
assign \phy_ddio_dqslogic_fiforeset[2]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[2];
assign \phy_ddio_dqslogic_fiforeset[3]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[3];

assign \phy_ddio_dqslogic_incrdataen[0]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[0];
assign \phy_ddio_dqslogic_incrdataen[1]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[1];
assign \phy_ddio_dqslogic_incrdataen[2]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[2];
assign \phy_ddio_dqslogic_incrdataen[3]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[3];
assign \phy_ddio_dqslogic_incrdataen[4]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[4];
assign \phy_ddio_dqslogic_incrdataen[5]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[5];
assign \phy_ddio_dqslogic_incrdataen[6]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[6];
assign \phy_ddio_dqslogic_incrdataen[7]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[7];

assign \phy_ddio_dqslogic_incwrptr[0]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[0];
assign \phy_ddio_dqslogic_incwrptr[1]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[1];
assign \phy_ddio_dqslogic_incwrptr[2]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[2];
assign \phy_ddio_dqslogic_incwrptr[3]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[3];
assign \phy_ddio_dqslogic_incwrptr[4]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[4];
assign \phy_ddio_dqslogic_incwrptr[5]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[5];
assign \phy_ddio_dqslogic_incwrptr[6]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[6];
assign \phy_ddio_dqslogic_incwrptr[7]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[7];

assign \phy_ddio_dqslogic_oct[0]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[0];
assign \phy_ddio_dqslogic_oct[1]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[1];
assign \phy_ddio_dqslogic_oct[2]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[2];
assign \phy_ddio_dqslogic_oct[3]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[3];
assign \phy_ddio_dqslogic_oct[4]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[4];
assign \phy_ddio_dqslogic_oct[5]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[5];
assign \phy_ddio_dqslogic_oct[6]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[6];
assign \phy_ddio_dqslogic_oct[7]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[7];

assign \phy_ddio_dqslogic_readlatency[0]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[0];
assign \phy_ddio_dqslogic_readlatency[1]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[1];
assign \phy_ddio_dqslogic_readlatency[2]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[2];
assign \phy_ddio_dqslogic_readlatency[3]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[3];
assign \phy_ddio_dqslogic_readlatency[4]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[4];
assign \phy_ddio_dqslogic_readlatency[5]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[5];
assign \phy_ddio_dqslogic_readlatency[6]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[6];
assign \phy_ddio_dqslogic_readlatency[7]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[7];
assign \phy_ddio_dqslogic_readlatency[8]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[8];
assign \phy_ddio_dqslogic_readlatency[9]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[9];
assign \phy_ddio_dqslogic_readlatency[10]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[10];
assign \phy_ddio_dqslogic_readlatency[11]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[11];
assign \phy_ddio_dqslogic_readlatency[12]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[12];
assign \phy_ddio_dqslogic_readlatency[13]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[13];
assign \phy_ddio_dqslogic_readlatency[14]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[14];
assign \phy_ddio_dqslogic_readlatency[15]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[15];
assign \phy_ddio_dqslogic_readlatency[16]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[16];
assign \phy_ddio_dqslogic_readlatency[17]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[17];
assign \phy_ddio_dqslogic_readlatency[18]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[18];
assign \phy_ddio_dqslogic_readlatency[19]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[19];

assign \phy_ddio_dqs_oe[0]  = hphy_inst_PHYDDIODQSOE_bus[0];
assign \phy_ddio_dqs_oe[1]  = hphy_inst_PHYDDIODQSOE_bus[1];
assign \phy_ddio_dqs_oe[2]  = hphy_inst_PHYDDIODQSOE_bus[2];
assign \phy_ddio_dqs_oe[3]  = hphy_inst_PHYDDIODQSOE_bus[3];
assign \phy_ddio_dqs_oe[4]  = hphy_inst_PHYDDIODQSOE_bus[4];
assign \phy_ddio_dqs_oe[5]  = hphy_inst_PHYDDIODQSOE_bus[5];
assign \phy_ddio_dqs_oe[6]  = hphy_inst_PHYDDIODQSOE_bus[6];
assign \phy_ddio_dqs_oe[7]  = hphy_inst_PHYDDIODQSOE_bus[7];

assign \phy_ddio_odt[0]  = hphy_inst_PHYDDIOODTDOUT_bus[0];
assign \phy_ddio_odt[1]  = hphy_inst_PHYDDIOODTDOUT_bus[1];
assign \phy_ddio_odt[2]  = hphy_inst_PHYDDIOODTDOUT_bus[2];
assign \phy_ddio_odt[3]  = hphy_inst_PHYDDIOODTDOUT_bus[3];

assign \phy_ddio_ras_n[0]  = hphy_inst_PHYDDIORASNDOUT_bus[0];
assign \phy_ddio_ras_n[1]  = hphy_inst_PHYDDIORASNDOUT_bus[1];
assign \phy_ddio_ras_n[2]  = hphy_inst_PHYDDIORASNDOUT_bus[2];
assign \phy_ddio_ras_n[3]  = hphy_inst_PHYDDIORASNDOUT_bus[3];

assign \phy_ddio_reset_n[0]  = hphy_inst_PHYDDIORESETNDOUT_bus[0];
assign \phy_ddio_reset_n[1]  = hphy_inst_PHYDDIORESETNDOUT_bus[1];
assign \phy_ddio_reset_n[2]  = hphy_inst_PHYDDIORESETNDOUT_bus[2];
assign \phy_ddio_reset_n[3]  = hphy_inst_PHYDDIORESETNDOUT_bus[3];

assign \phy_ddio_we_n[0]  = hphy_inst_PHYDDIOWENDOUT_bus[0];
assign \phy_ddio_we_n[1]  = hphy_inst_PHYDDIOWENDOUT_bus[1];
assign \phy_ddio_we_n[2]  = hphy_inst_PHYDDIOWENDOUT_bus[2];
assign \phy_ddio_we_n[3]  = hphy_inst_PHYDDIOWENDOUT_bus[3];

system_hps_sdram_p0_acv_hard_io_pads uio_pads(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(\phy_ddio_address[0] ),
	.phy_ddio_address_1(\phy_ddio_address[1] ),
	.phy_ddio_address_2(\phy_ddio_address[2] ),
	.phy_ddio_address_3(\phy_ddio_address[3] ),
	.phy_ddio_address_4(\phy_ddio_address[4] ),
	.phy_ddio_address_5(\phy_ddio_address[5] ),
	.phy_ddio_address_6(\phy_ddio_address[6] ),
	.phy_ddio_address_7(\phy_ddio_address[7] ),
	.phy_ddio_address_8(\phy_ddio_address[8] ),
	.phy_ddio_address_9(\phy_ddio_address[9] ),
	.phy_ddio_address_10(\phy_ddio_address[10] ),
	.phy_ddio_address_11(\phy_ddio_address[11] ),
	.phy_ddio_address_12(\phy_ddio_address[12] ),
	.phy_ddio_address_13(\phy_ddio_address[13] ),
	.phy_ddio_address_14(\phy_ddio_address[14] ),
	.phy_ddio_address_15(\phy_ddio_address[15] ),
	.phy_ddio_address_16(\phy_ddio_address[16] ),
	.phy_ddio_address_17(\phy_ddio_address[17] ),
	.phy_ddio_address_18(\phy_ddio_address[18] ),
	.phy_ddio_address_19(\phy_ddio_address[19] ),
	.phy_ddio_address_20(\phy_ddio_address[20] ),
	.phy_ddio_address_21(\phy_ddio_address[21] ),
	.phy_ddio_address_22(\phy_ddio_address[22] ),
	.phy_ddio_address_23(\phy_ddio_address[23] ),
	.phy_ddio_address_24(\phy_ddio_address[24] ),
	.phy_ddio_address_25(\phy_ddio_address[25] ),
	.phy_ddio_address_26(\phy_ddio_address[26] ),
	.phy_ddio_address_27(\phy_ddio_address[27] ),
	.phy_ddio_address_28(\phy_ddio_address[28] ),
	.phy_ddio_address_29(\phy_ddio_address[29] ),
	.phy_ddio_address_30(\phy_ddio_address[30] ),
	.phy_ddio_address_31(\phy_ddio_address[31] ),
	.phy_ddio_address_32(\phy_ddio_address[32] ),
	.phy_ddio_address_33(\phy_ddio_address[33] ),
	.phy_ddio_address_34(\phy_ddio_address[34] ),
	.phy_ddio_address_35(\phy_ddio_address[35] ),
	.phy_ddio_address_36(\phy_ddio_address[36] ),
	.phy_ddio_address_37(\phy_ddio_address[37] ),
	.phy_ddio_address_38(\phy_ddio_address[38] ),
	.phy_ddio_address_39(\phy_ddio_address[39] ),
	.phy_ddio_address_40(\phy_ddio_address[40] ),
	.phy_ddio_address_41(\phy_ddio_address[41] ),
	.phy_ddio_address_42(\phy_ddio_address[42] ),
	.phy_ddio_address_43(\phy_ddio_address[43] ),
	.phy_ddio_address_44(\phy_ddio_address[44] ),
	.phy_ddio_address_45(\phy_ddio_address[45] ),
	.phy_ddio_address_46(\phy_ddio_address[46] ),
	.phy_ddio_address_47(\phy_ddio_address[47] ),
	.phy_ddio_address_48(\phy_ddio_address[48] ),
	.phy_ddio_address_49(\phy_ddio_address[49] ),
	.phy_ddio_address_50(\phy_ddio_address[50] ),
	.phy_ddio_address_51(\phy_ddio_address[51] ),
	.phy_ddio_address_52(\phy_ddio_address[52] ),
	.phy_ddio_address_53(\phy_ddio_address[53] ),
	.phy_ddio_address_54(\phy_ddio_address[54] ),
	.phy_ddio_address_55(\phy_ddio_address[55] ),
	.phy_ddio_address_56(\phy_ddio_address[56] ),
	.phy_ddio_address_57(\phy_ddio_address[57] ),
	.phy_ddio_address_58(\phy_ddio_address[58] ),
	.phy_ddio_address_59(\phy_ddio_address[59] ),
	.phy_ddio_bank_0(\phy_ddio_bank[0] ),
	.phy_ddio_bank_1(\phy_ddio_bank[1] ),
	.phy_ddio_bank_2(\phy_ddio_bank[2] ),
	.phy_ddio_bank_3(\phy_ddio_bank[3] ),
	.phy_ddio_bank_4(\phy_ddio_bank[4] ),
	.phy_ddio_bank_5(\phy_ddio_bank[5] ),
	.phy_ddio_bank_6(\phy_ddio_bank[6] ),
	.phy_ddio_bank_7(\phy_ddio_bank[7] ),
	.phy_ddio_bank_8(\phy_ddio_bank[8] ),
	.phy_ddio_bank_9(\phy_ddio_bank[9] ),
	.phy_ddio_bank_10(\phy_ddio_bank[10] ),
	.phy_ddio_bank_11(\phy_ddio_bank[11] ),
	.phy_ddio_cas_n_0(\phy_ddio_cas_n[0] ),
	.phy_ddio_cas_n_1(\phy_ddio_cas_n[1] ),
	.phy_ddio_cas_n_2(\phy_ddio_cas_n[2] ),
	.phy_ddio_cas_n_3(\phy_ddio_cas_n[3] ),
	.phy_ddio_ck_0(\phy_ddio_ck[0] ),
	.phy_ddio_ck_1(\phy_ddio_ck[1] ),
	.phy_ddio_cke_0(\phy_ddio_cke[0] ),
	.phy_ddio_cke_1(\phy_ddio_cke[1] ),
	.phy_ddio_cke_2(\phy_ddio_cke[2] ),
	.phy_ddio_cke_3(\phy_ddio_cke[3] ),
	.phy_ddio_cs_n_0(\phy_ddio_cs_n[0] ),
	.phy_ddio_cs_n_1(\phy_ddio_cs_n[1] ),
	.phy_ddio_cs_n_2(\phy_ddio_cs_n[2] ),
	.phy_ddio_cs_n_3(\phy_ddio_cs_n[3] ),
	.phy_ddio_dmdout_0(\phy_ddio_dmdout[0] ),
	.phy_ddio_dmdout_1(\phy_ddio_dmdout[1] ),
	.phy_ddio_dmdout_2(\phy_ddio_dmdout[2] ),
	.phy_ddio_dmdout_3(\phy_ddio_dmdout[3] ),
	.phy_ddio_dmdout_4(\phy_ddio_dmdout[4] ),
	.phy_ddio_dmdout_5(\phy_ddio_dmdout[5] ),
	.phy_ddio_dmdout_6(\phy_ddio_dmdout[6] ),
	.phy_ddio_dmdout_7(\phy_ddio_dmdout[7] ),
	.phy_ddio_dmdout_8(\phy_ddio_dmdout[8] ),
	.phy_ddio_dmdout_9(\phy_ddio_dmdout[9] ),
	.phy_ddio_dmdout_10(\phy_ddio_dmdout[10] ),
	.phy_ddio_dmdout_11(\phy_ddio_dmdout[11] ),
	.phy_ddio_dmdout_12(\phy_ddio_dmdout[12] ),
	.phy_ddio_dmdout_13(\phy_ddio_dmdout[13] ),
	.phy_ddio_dmdout_14(\phy_ddio_dmdout[14] ),
	.phy_ddio_dmdout_15(\phy_ddio_dmdout[15] ),
	.phy_ddio_dqdout_0(\phy_ddio_dqdout[0] ),
	.phy_ddio_dqdout_1(\phy_ddio_dqdout[1] ),
	.phy_ddio_dqdout_2(\phy_ddio_dqdout[2] ),
	.phy_ddio_dqdout_3(\phy_ddio_dqdout[3] ),
	.phy_ddio_dqdout_4(\phy_ddio_dqdout[4] ),
	.phy_ddio_dqdout_5(\phy_ddio_dqdout[5] ),
	.phy_ddio_dqdout_6(\phy_ddio_dqdout[6] ),
	.phy_ddio_dqdout_7(\phy_ddio_dqdout[7] ),
	.phy_ddio_dqdout_8(\phy_ddio_dqdout[8] ),
	.phy_ddio_dqdout_9(\phy_ddio_dqdout[9] ),
	.phy_ddio_dqdout_10(\phy_ddio_dqdout[10] ),
	.phy_ddio_dqdout_11(\phy_ddio_dqdout[11] ),
	.phy_ddio_dqdout_12(\phy_ddio_dqdout[12] ),
	.phy_ddio_dqdout_13(\phy_ddio_dqdout[13] ),
	.phy_ddio_dqdout_14(\phy_ddio_dqdout[14] ),
	.phy_ddio_dqdout_15(\phy_ddio_dqdout[15] ),
	.phy_ddio_dqdout_16(\phy_ddio_dqdout[16] ),
	.phy_ddio_dqdout_17(\phy_ddio_dqdout[17] ),
	.phy_ddio_dqdout_18(\phy_ddio_dqdout[18] ),
	.phy_ddio_dqdout_19(\phy_ddio_dqdout[19] ),
	.phy_ddio_dqdout_20(\phy_ddio_dqdout[20] ),
	.phy_ddio_dqdout_21(\phy_ddio_dqdout[21] ),
	.phy_ddio_dqdout_22(\phy_ddio_dqdout[22] ),
	.phy_ddio_dqdout_23(\phy_ddio_dqdout[23] ),
	.phy_ddio_dqdout_24(\phy_ddio_dqdout[24] ),
	.phy_ddio_dqdout_25(\phy_ddio_dqdout[25] ),
	.phy_ddio_dqdout_26(\phy_ddio_dqdout[26] ),
	.phy_ddio_dqdout_27(\phy_ddio_dqdout[27] ),
	.phy_ddio_dqdout_28(\phy_ddio_dqdout[28] ),
	.phy_ddio_dqdout_29(\phy_ddio_dqdout[29] ),
	.phy_ddio_dqdout_30(\phy_ddio_dqdout[30] ),
	.phy_ddio_dqdout_31(\phy_ddio_dqdout[31] ),
	.phy_ddio_dqdout_36(\phy_ddio_dqdout[36] ),
	.phy_ddio_dqdout_37(\phy_ddio_dqdout[37] ),
	.phy_ddio_dqdout_38(\phy_ddio_dqdout[38] ),
	.phy_ddio_dqdout_39(\phy_ddio_dqdout[39] ),
	.phy_ddio_dqdout_40(\phy_ddio_dqdout[40] ),
	.phy_ddio_dqdout_41(\phy_ddio_dqdout[41] ),
	.phy_ddio_dqdout_42(\phy_ddio_dqdout[42] ),
	.phy_ddio_dqdout_43(\phy_ddio_dqdout[43] ),
	.phy_ddio_dqdout_44(\phy_ddio_dqdout[44] ),
	.phy_ddio_dqdout_45(\phy_ddio_dqdout[45] ),
	.phy_ddio_dqdout_46(\phy_ddio_dqdout[46] ),
	.phy_ddio_dqdout_47(\phy_ddio_dqdout[47] ),
	.phy_ddio_dqdout_48(\phy_ddio_dqdout[48] ),
	.phy_ddio_dqdout_49(\phy_ddio_dqdout[49] ),
	.phy_ddio_dqdout_50(\phy_ddio_dqdout[50] ),
	.phy_ddio_dqdout_51(\phy_ddio_dqdout[51] ),
	.phy_ddio_dqdout_52(\phy_ddio_dqdout[52] ),
	.phy_ddio_dqdout_53(\phy_ddio_dqdout[53] ),
	.phy_ddio_dqdout_54(\phy_ddio_dqdout[54] ),
	.phy_ddio_dqdout_55(\phy_ddio_dqdout[55] ),
	.phy_ddio_dqdout_56(\phy_ddio_dqdout[56] ),
	.phy_ddio_dqdout_57(\phy_ddio_dqdout[57] ),
	.phy_ddio_dqdout_58(\phy_ddio_dqdout[58] ),
	.phy_ddio_dqdout_59(\phy_ddio_dqdout[59] ),
	.phy_ddio_dqdout_60(\phy_ddio_dqdout[60] ),
	.phy_ddio_dqdout_61(\phy_ddio_dqdout[61] ),
	.phy_ddio_dqdout_62(\phy_ddio_dqdout[62] ),
	.phy_ddio_dqdout_63(\phy_ddio_dqdout[63] ),
	.phy_ddio_dqdout_64(\phy_ddio_dqdout[64] ),
	.phy_ddio_dqdout_65(\phy_ddio_dqdout[65] ),
	.phy_ddio_dqdout_66(\phy_ddio_dqdout[66] ),
	.phy_ddio_dqdout_67(\phy_ddio_dqdout[67] ),
	.phy_ddio_dqdout_72(\phy_ddio_dqdout[72] ),
	.phy_ddio_dqdout_73(\phy_ddio_dqdout[73] ),
	.phy_ddio_dqdout_74(\phy_ddio_dqdout[74] ),
	.phy_ddio_dqdout_75(\phy_ddio_dqdout[75] ),
	.phy_ddio_dqdout_76(\phy_ddio_dqdout[76] ),
	.phy_ddio_dqdout_77(\phy_ddio_dqdout[77] ),
	.phy_ddio_dqdout_78(\phy_ddio_dqdout[78] ),
	.phy_ddio_dqdout_79(\phy_ddio_dqdout[79] ),
	.phy_ddio_dqdout_80(\phy_ddio_dqdout[80] ),
	.phy_ddio_dqdout_81(\phy_ddio_dqdout[81] ),
	.phy_ddio_dqdout_82(\phy_ddio_dqdout[82] ),
	.phy_ddio_dqdout_83(\phy_ddio_dqdout[83] ),
	.phy_ddio_dqdout_84(\phy_ddio_dqdout[84] ),
	.phy_ddio_dqdout_85(\phy_ddio_dqdout[85] ),
	.phy_ddio_dqdout_86(\phy_ddio_dqdout[86] ),
	.phy_ddio_dqdout_87(\phy_ddio_dqdout[87] ),
	.phy_ddio_dqdout_88(\phy_ddio_dqdout[88] ),
	.phy_ddio_dqdout_89(\phy_ddio_dqdout[89] ),
	.phy_ddio_dqdout_90(\phy_ddio_dqdout[90] ),
	.phy_ddio_dqdout_91(\phy_ddio_dqdout[91] ),
	.phy_ddio_dqdout_92(\phy_ddio_dqdout[92] ),
	.phy_ddio_dqdout_93(\phy_ddio_dqdout[93] ),
	.phy_ddio_dqdout_94(\phy_ddio_dqdout[94] ),
	.phy_ddio_dqdout_95(\phy_ddio_dqdout[95] ),
	.phy_ddio_dqdout_96(\phy_ddio_dqdout[96] ),
	.phy_ddio_dqdout_97(\phy_ddio_dqdout[97] ),
	.phy_ddio_dqdout_98(\phy_ddio_dqdout[98] ),
	.phy_ddio_dqdout_99(\phy_ddio_dqdout[99] ),
	.phy_ddio_dqdout_100(\phy_ddio_dqdout[100] ),
	.phy_ddio_dqdout_101(\phy_ddio_dqdout[101] ),
	.phy_ddio_dqdout_102(\phy_ddio_dqdout[102] ),
	.phy_ddio_dqdout_103(\phy_ddio_dqdout[103] ),
	.phy_ddio_dqdout_108(\phy_ddio_dqdout[108] ),
	.phy_ddio_dqdout_109(\phy_ddio_dqdout[109] ),
	.phy_ddio_dqdout_110(\phy_ddio_dqdout[110] ),
	.phy_ddio_dqdout_111(\phy_ddio_dqdout[111] ),
	.phy_ddio_dqdout_112(\phy_ddio_dqdout[112] ),
	.phy_ddio_dqdout_113(\phy_ddio_dqdout[113] ),
	.phy_ddio_dqdout_114(\phy_ddio_dqdout[114] ),
	.phy_ddio_dqdout_115(\phy_ddio_dqdout[115] ),
	.phy_ddio_dqdout_116(\phy_ddio_dqdout[116] ),
	.phy_ddio_dqdout_117(\phy_ddio_dqdout[117] ),
	.phy_ddio_dqdout_118(\phy_ddio_dqdout[118] ),
	.phy_ddio_dqdout_119(\phy_ddio_dqdout[119] ),
	.phy_ddio_dqdout_120(\phy_ddio_dqdout[120] ),
	.phy_ddio_dqdout_121(\phy_ddio_dqdout[121] ),
	.phy_ddio_dqdout_122(\phy_ddio_dqdout[122] ),
	.phy_ddio_dqdout_123(\phy_ddio_dqdout[123] ),
	.phy_ddio_dqdout_124(\phy_ddio_dqdout[124] ),
	.phy_ddio_dqdout_125(\phy_ddio_dqdout[125] ),
	.phy_ddio_dqdout_126(\phy_ddio_dqdout[126] ),
	.phy_ddio_dqdout_127(\phy_ddio_dqdout[127] ),
	.phy_ddio_dqdout_128(\phy_ddio_dqdout[128] ),
	.phy_ddio_dqdout_129(\phy_ddio_dqdout[129] ),
	.phy_ddio_dqdout_130(\phy_ddio_dqdout[130] ),
	.phy_ddio_dqdout_131(\phy_ddio_dqdout[131] ),
	.phy_ddio_dqdout_132(\phy_ddio_dqdout[132] ),
	.phy_ddio_dqdout_133(\phy_ddio_dqdout[133] ),
	.phy_ddio_dqdout_134(\phy_ddio_dqdout[134] ),
	.phy_ddio_dqdout_135(\phy_ddio_dqdout[135] ),
	.phy_ddio_dqdout_136(\phy_ddio_dqdout[136] ),
	.phy_ddio_dqdout_137(\phy_ddio_dqdout[137] ),
	.phy_ddio_dqdout_138(\phy_ddio_dqdout[138] ),
	.phy_ddio_dqdout_139(\phy_ddio_dqdout[139] ),
	.phy_ddio_dqoe_0(\phy_ddio_dqoe[0] ),
	.phy_ddio_dqoe_1(\phy_ddio_dqoe[1] ),
	.phy_ddio_dqoe_2(\phy_ddio_dqoe[2] ),
	.phy_ddio_dqoe_3(\phy_ddio_dqoe[3] ),
	.phy_ddio_dqoe_4(\phy_ddio_dqoe[4] ),
	.phy_ddio_dqoe_5(\phy_ddio_dqoe[5] ),
	.phy_ddio_dqoe_6(\phy_ddio_dqoe[6] ),
	.phy_ddio_dqoe_7(\phy_ddio_dqoe[7] ),
	.phy_ddio_dqoe_8(\phy_ddio_dqoe[8] ),
	.phy_ddio_dqoe_9(\phy_ddio_dqoe[9] ),
	.phy_ddio_dqoe_10(\phy_ddio_dqoe[10] ),
	.phy_ddio_dqoe_11(\phy_ddio_dqoe[11] ),
	.phy_ddio_dqoe_12(\phy_ddio_dqoe[12] ),
	.phy_ddio_dqoe_13(\phy_ddio_dqoe[13] ),
	.phy_ddio_dqoe_14(\phy_ddio_dqoe[14] ),
	.phy_ddio_dqoe_15(\phy_ddio_dqoe[15] ),
	.phy_ddio_dqoe_18(\phy_ddio_dqoe[18] ),
	.phy_ddio_dqoe_19(\phy_ddio_dqoe[19] ),
	.phy_ddio_dqoe_20(\phy_ddio_dqoe[20] ),
	.phy_ddio_dqoe_21(\phy_ddio_dqoe[21] ),
	.phy_ddio_dqoe_22(\phy_ddio_dqoe[22] ),
	.phy_ddio_dqoe_23(\phy_ddio_dqoe[23] ),
	.phy_ddio_dqoe_24(\phy_ddio_dqoe[24] ),
	.phy_ddio_dqoe_25(\phy_ddio_dqoe[25] ),
	.phy_ddio_dqoe_26(\phy_ddio_dqoe[26] ),
	.phy_ddio_dqoe_27(\phy_ddio_dqoe[27] ),
	.phy_ddio_dqoe_28(\phy_ddio_dqoe[28] ),
	.phy_ddio_dqoe_29(\phy_ddio_dqoe[29] ),
	.phy_ddio_dqoe_30(\phy_ddio_dqoe[30] ),
	.phy_ddio_dqoe_31(\phy_ddio_dqoe[31] ),
	.phy_ddio_dqoe_32(\phy_ddio_dqoe[32] ),
	.phy_ddio_dqoe_33(\phy_ddio_dqoe[33] ),
	.phy_ddio_dqoe_36(\phy_ddio_dqoe[36] ),
	.phy_ddio_dqoe_37(\phy_ddio_dqoe[37] ),
	.phy_ddio_dqoe_38(\phy_ddio_dqoe[38] ),
	.phy_ddio_dqoe_39(\phy_ddio_dqoe[39] ),
	.phy_ddio_dqoe_40(\phy_ddio_dqoe[40] ),
	.phy_ddio_dqoe_41(\phy_ddio_dqoe[41] ),
	.phy_ddio_dqoe_42(\phy_ddio_dqoe[42] ),
	.phy_ddio_dqoe_43(\phy_ddio_dqoe[43] ),
	.phy_ddio_dqoe_44(\phy_ddio_dqoe[44] ),
	.phy_ddio_dqoe_45(\phy_ddio_dqoe[45] ),
	.phy_ddio_dqoe_46(\phy_ddio_dqoe[46] ),
	.phy_ddio_dqoe_47(\phy_ddio_dqoe[47] ),
	.phy_ddio_dqoe_48(\phy_ddio_dqoe[48] ),
	.phy_ddio_dqoe_49(\phy_ddio_dqoe[49] ),
	.phy_ddio_dqoe_50(\phy_ddio_dqoe[50] ),
	.phy_ddio_dqoe_51(\phy_ddio_dqoe[51] ),
	.phy_ddio_dqoe_54(\phy_ddio_dqoe[54] ),
	.phy_ddio_dqoe_55(\phy_ddio_dqoe[55] ),
	.phy_ddio_dqoe_56(\phy_ddio_dqoe[56] ),
	.phy_ddio_dqoe_57(\phy_ddio_dqoe[57] ),
	.phy_ddio_dqoe_58(\phy_ddio_dqoe[58] ),
	.phy_ddio_dqoe_59(\phy_ddio_dqoe[59] ),
	.phy_ddio_dqoe_60(\phy_ddio_dqoe[60] ),
	.phy_ddio_dqoe_61(\phy_ddio_dqoe[61] ),
	.phy_ddio_dqoe_62(\phy_ddio_dqoe[62] ),
	.phy_ddio_dqoe_63(\phy_ddio_dqoe[63] ),
	.phy_ddio_dqoe_64(\phy_ddio_dqoe[64] ),
	.phy_ddio_dqoe_65(\phy_ddio_dqoe[65] ),
	.phy_ddio_dqoe_66(\phy_ddio_dqoe[66] ),
	.phy_ddio_dqoe_67(\phy_ddio_dqoe[67] ),
	.phy_ddio_dqoe_68(\phy_ddio_dqoe[68] ),
	.phy_ddio_dqoe_69(\phy_ddio_dqoe[69] ),
	.phy_ddio_dqs_dout_0(\phy_ddio_dqs_dout[0] ),
	.phy_ddio_dqs_dout_1(\phy_ddio_dqs_dout[1] ),
	.phy_ddio_dqs_dout_2(\phy_ddio_dqs_dout[2] ),
	.phy_ddio_dqs_dout_3(\phy_ddio_dqs_dout[3] ),
	.phy_ddio_dqs_dout_4(\phy_ddio_dqs_dout[4] ),
	.phy_ddio_dqs_dout_5(\phy_ddio_dqs_dout[5] ),
	.phy_ddio_dqs_dout_6(\phy_ddio_dqs_dout[6] ),
	.phy_ddio_dqs_dout_7(\phy_ddio_dqs_dout[7] ),
	.phy_ddio_dqs_dout_8(\phy_ddio_dqs_dout[8] ),
	.phy_ddio_dqs_dout_9(\phy_ddio_dqs_dout[9] ),
	.phy_ddio_dqs_dout_10(\phy_ddio_dqs_dout[10] ),
	.phy_ddio_dqs_dout_11(\phy_ddio_dqs_dout[11] ),
	.phy_ddio_dqs_dout_12(\phy_ddio_dqs_dout[12] ),
	.phy_ddio_dqs_dout_13(\phy_ddio_dqs_dout[13] ),
	.phy_ddio_dqs_dout_14(\phy_ddio_dqs_dout[14] ),
	.phy_ddio_dqs_dout_15(\phy_ddio_dqs_dout[15] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(\phy_ddio_dqslogic_aclr_fifoctrl[0] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(\phy_ddio_dqslogic_aclr_fifoctrl[1] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(\phy_ddio_dqslogic_aclr_fifoctrl[2] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(\phy_ddio_dqslogic_aclr_fifoctrl[3] ),
	.phy_ddio_dqslogic_aclr_pstamble_0(\phy_ddio_dqslogic_aclr_pstamble[0] ),
	.phy_ddio_dqslogic_aclr_pstamble_1(\phy_ddio_dqslogic_aclr_pstamble[1] ),
	.phy_ddio_dqslogic_aclr_pstamble_2(\phy_ddio_dqslogic_aclr_pstamble[2] ),
	.phy_ddio_dqslogic_aclr_pstamble_3(\phy_ddio_dqslogic_aclr_pstamble[3] ),
	.phy_ddio_dqslogic_dqsena_0(\phy_ddio_dqslogic_dqsena[0] ),
	.phy_ddio_dqslogic_dqsena_1(\phy_ddio_dqslogic_dqsena[1] ),
	.phy_ddio_dqslogic_dqsena_2(\phy_ddio_dqslogic_dqsena[2] ),
	.phy_ddio_dqslogic_dqsena_3(\phy_ddio_dqslogic_dqsena[3] ),
	.phy_ddio_dqslogic_dqsena_4(\phy_ddio_dqslogic_dqsena[4] ),
	.phy_ddio_dqslogic_dqsena_5(\phy_ddio_dqslogic_dqsena[5] ),
	.phy_ddio_dqslogic_dqsena_6(\phy_ddio_dqslogic_dqsena[6] ),
	.phy_ddio_dqslogic_dqsena_7(\phy_ddio_dqslogic_dqsena[7] ),
	.phy_ddio_dqslogic_fiforeset_0(\phy_ddio_dqslogic_fiforeset[0] ),
	.phy_ddio_dqslogic_fiforeset_1(\phy_ddio_dqslogic_fiforeset[1] ),
	.phy_ddio_dqslogic_fiforeset_2(\phy_ddio_dqslogic_fiforeset[2] ),
	.phy_ddio_dqslogic_fiforeset_3(\phy_ddio_dqslogic_fiforeset[3] ),
	.phy_ddio_dqslogic_incrdataen_0(\phy_ddio_dqslogic_incrdataen[0] ),
	.phy_ddio_dqslogic_incrdataen_1(\phy_ddio_dqslogic_incrdataen[1] ),
	.phy_ddio_dqslogic_incrdataen_2(\phy_ddio_dqslogic_incrdataen[2] ),
	.phy_ddio_dqslogic_incrdataen_3(\phy_ddio_dqslogic_incrdataen[3] ),
	.phy_ddio_dqslogic_incrdataen_4(\phy_ddio_dqslogic_incrdataen[4] ),
	.phy_ddio_dqslogic_incrdataen_5(\phy_ddio_dqslogic_incrdataen[5] ),
	.phy_ddio_dqslogic_incrdataen_6(\phy_ddio_dqslogic_incrdataen[6] ),
	.phy_ddio_dqslogic_incrdataen_7(\phy_ddio_dqslogic_incrdataen[7] ),
	.phy_ddio_dqslogic_incwrptr_0(\phy_ddio_dqslogic_incwrptr[0] ),
	.phy_ddio_dqslogic_incwrptr_1(\phy_ddio_dqslogic_incwrptr[1] ),
	.phy_ddio_dqslogic_incwrptr_2(\phy_ddio_dqslogic_incwrptr[2] ),
	.phy_ddio_dqslogic_incwrptr_3(\phy_ddio_dqslogic_incwrptr[3] ),
	.phy_ddio_dqslogic_incwrptr_4(\phy_ddio_dqslogic_incwrptr[4] ),
	.phy_ddio_dqslogic_incwrptr_5(\phy_ddio_dqslogic_incwrptr[5] ),
	.phy_ddio_dqslogic_incwrptr_6(\phy_ddio_dqslogic_incwrptr[6] ),
	.phy_ddio_dqslogic_incwrptr_7(\phy_ddio_dqslogic_incwrptr[7] ),
	.phy_ddio_dqslogic_oct_0(\phy_ddio_dqslogic_oct[0] ),
	.phy_ddio_dqslogic_oct_1(\phy_ddio_dqslogic_oct[1] ),
	.phy_ddio_dqslogic_oct_2(\phy_ddio_dqslogic_oct[2] ),
	.phy_ddio_dqslogic_oct_3(\phy_ddio_dqslogic_oct[3] ),
	.phy_ddio_dqslogic_oct_4(\phy_ddio_dqslogic_oct[4] ),
	.phy_ddio_dqslogic_oct_5(\phy_ddio_dqslogic_oct[5] ),
	.phy_ddio_dqslogic_oct_6(\phy_ddio_dqslogic_oct[6] ),
	.phy_ddio_dqslogic_oct_7(\phy_ddio_dqslogic_oct[7] ),
	.phy_ddio_dqslogic_readlatency_0(\phy_ddio_dqslogic_readlatency[0] ),
	.phy_ddio_dqslogic_readlatency_1(\phy_ddio_dqslogic_readlatency[1] ),
	.phy_ddio_dqslogic_readlatency_2(\phy_ddio_dqslogic_readlatency[2] ),
	.phy_ddio_dqslogic_readlatency_3(\phy_ddio_dqslogic_readlatency[3] ),
	.phy_ddio_dqslogic_readlatency_4(\phy_ddio_dqslogic_readlatency[4] ),
	.phy_ddio_dqslogic_readlatency_5(\phy_ddio_dqslogic_readlatency[5] ),
	.phy_ddio_dqslogic_readlatency_6(\phy_ddio_dqslogic_readlatency[6] ),
	.phy_ddio_dqslogic_readlatency_7(\phy_ddio_dqslogic_readlatency[7] ),
	.phy_ddio_dqslogic_readlatency_8(\phy_ddio_dqslogic_readlatency[8] ),
	.phy_ddio_dqslogic_readlatency_9(\phy_ddio_dqslogic_readlatency[9] ),
	.phy_ddio_dqslogic_readlatency_10(\phy_ddio_dqslogic_readlatency[10] ),
	.phy_ddio_dqslogic_readlatency_11(\phy_ddio_dqslogic_readlatency[11] ),
	.phy_ddio_dqslogic_readlatency_12(\phy_ddio_dqslogic_readlatency[12] ),
	.phy_ddio_dqslogic_readlatency_13(\phy_ddio_dqslogic_readlatency[13] ),
	.phy_ddio_dqslogic_readlatency_14(\phy_ddio_dqslogic_readlatency[14] ),
	.phy_ddio_dqslogic_readlatency_15(\phy_ddio_dqslogic_readlatency[15] ),
	.phy_ddio_dqslogic_readlatency_16(\phy_ddio_dqslogic_readlatency[16] ),
	.phy_ddio_dqslogic_readlatency_17(\phy_ddio_dqslogic_readlatency[17] ),
	.phy_ddio_dqslogic_readlatency_18(\phy_ddio_dqslogic_readlatency[18] ),
	.phy_ddio_dqslogic_readlatency_19(\phy_ddio_dqslogic_readlatency[19] ),
	.phy_ddio_dqs_oe_0(\phy_ddio_dqs_oe[0] ),
	.phy_ddio_dqs_oe_1(\phy_ddio_dqs_oe[1] ),
	.phy_ddio_dqs_oe_2(\phy_ddio_dqs_oe[2] ),
	.phy_ddio_dqs_oe_3(\phy_ddio_dqs_oe[3] ),
	.phy_ddio_dqs_oe_4(\phy_ddio_dqs_oe[4] ),
	.phy_ddio_dqs_oe_5(\phy_ddio_dqs_oe[5] ),
	.phy_ddio_dqs_oe_6(\phy_ddio_dqs_oe[6] ),
	.phy_ddio_dqs_oe_7(\phy_ddio_dqs_oe[7] ),
	.phy_ddio_odt_0(\phy_ddio_odt[0] ),
	.phy_ddio_odt_1(\phy_ddio_odt[1] ),
	.phy_ddio_odt_2(\phy_ddio_odt[2] ),
	.phy_ddio_odt_3(\phy_ddio_odt[3] ),
	.phy_ddio_ras_n_0(\phy_ddio_ras_n[0] ),
	.phy_ddio_ras_n_1(\phy_ddio_ras_n[1] ),
	.phy_ddio_ras_n_2(\phy_ddio_ras_n[2] ),
	.phy_ddio_ras_n_3(\phy_ddio_ras_n[3] ),
	.phy_ddio_reset_n_0(\phy_ddio_reset_n[0] ),
	.phy_ddio_reset_n_1(\phy_ddio_reset_n[1] ),
	.phy_ddio_reset_n_2(\phy_ddio_reset_n[2] ),
	.phy_ddio_reset_n_3(\phy_ddio_reset_n[3] ),
	.phy_ddio_we_n_0(\phy_ddio_we_n[0] ),
	.phy_ddio_we_n_1(\phy_ddio_we_n[1] ),
	.phy_ddio_we_n_2(\phy_ddio_we_n[2] ),
	.phy_ddio_we_n_3(\phy_ddio_we_n[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.ddio_phy_dqslogic_rdatavalid({ddio_phy_dqslogic_rdatavalid_unconnected_wire_4,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

system_hps_sdram_p0_acv_ldc_25 memphy_ldc(
	.pll_hr_clk(afi_clk),
	.pll_dqs_clk(afi_clk),
	.adc_clk(leveled_dqs_clocks_0),
	.avl_clk(\memphy_ldc|leveled_hr_clocks[0] ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_mem_phy hphy_inst(
	.aficasn(afi_cas_n[0]),
	.afimemclkdisable(afi_mem_clk_disable[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.avlread(gnd),
	.avlresetn(gnd),
	.avlwrite(gnd),
	.globalresetn(gnd),
	.iointcasnaclr(gnd),
	.iointrasnaclr(gnd),
	.iointresetnaclr(gnd),
	.iointwenaclr(gnd),
	.plladdrcmdclk(!leveled_dqs_clocks_0),
	.pllaficlk(leveled_dqs_clocks_0),
	.pllavlclk(\memphy_ldc|leveled_hr_clocks[0] ),
	.plllocked(gnd),
	.scanen(gnd),
	.softresetn(gnd),
	.afiaddr({afi_addr[19],afi_addr[18],afi_addr[17],afi_addr[16],afi_addr[15],afi_addr[14],afi_addr[13],afi_addr[12],afi_addr[11],afi_addr[10],afi_addr[9],afi_addr[8],afi_addr[7],afi_addr[6],afi_addr[5],afi_addr[4],afi_addr[3],afi_addr[2],afi_addr[1],afi_addr[0]}),
	.afiba({afi_ba[2],afi_ba[1],afi_ba[0]}),
	.aficke({afi_cke[1],afi_cke[0]}),
	.aficsn({afi_cs_n[1],afi_cs_n[0]}),
	.afidm({afi_dm[9],afi_dm[8],afi_dm[7],afi_dm[6],afi_dm[5],afi_dm[4],afi_dm[3],afi_dm[2],afi_dm[1],afi_dm[0]}),
	.afidqsburst({afi_dqs_burst[4],afi_dqs_burst[3],afi_dqs_burst[2],afi_dqs_burst[1],afi_dqs_burst[0]}),
	.afiodt({afi_odt[1],afi_odt[0]}),
	.afirdataen({afi_rdata_en[4],afi_rdata_en[3],afi_rdata_en[2],afi_rdata_en[1],afi_rdata_en[0]}),
	.afirdataenfull({afi_rdata_en_full[4],afi_rdata_en_full[3],afi_rdata_en_full[2],afi_rdata_en_full[1],afi_rdata_en_full[0]}),
	.afiwdata({afi_wdata[79],afi_wdata[78],afi_wdata[77],afi_wdata[76],afi_wdata[75],afi_wdata[74],afi_wdata[73],afi_wdata[72],afi_wdata[71],afi_wdata[70],afi_wdata[69],afi_wdata[68],afi_wdata[67],afi_wdata[66],afi_wdata[65],afi_wdata[64],afi_wdata[63],afi_wdata[62],afi_wdata[61],afi_wdata[60],afi_wdata[59],afi_wdata[58],afi_wdata[57],afi_wdata[56],afi_wdata[55],afi_wdata[54],afi_wdata[53],afi_wdata[52],
afi_wdata[51],afi_wdata[50],afi_wdata[49],afi_wdata[48],afi_wdata[47],afi_wdata[46],afi_wdata[45],afi_wdata[44],afi_wdata[43],afi_wdata[42],afi_wdata[41],afi_wdata[40],afi_wdata[39],afi_wdata[38],afi_wdata[37],afi_wdata[36],afi_wdata[35],afi_wdata[34],afi_wdata[33],afi_wdata[32],afi_wdata[31],afi_wdata[30],afi_wdata[29],afi_wdata[28],afi_wdata[27],afi_wdata[26],afi_wdata[25],afi_wdata[24],
afi_wdata[23],afi_wdata[22],afi_wdata[21],afi_wdata[20],afi_wdata[19],afi_wdata[18],afi_wdata[17],afi_wdata[16],afi_wdata[15],afi_wdata[14],afi_wdata[13],afi_wdata[12],afi_wdata[11],afi_wdata[10],afi_wdata[9],afi_wdata[8],afi_wdata[7],afi_wdata[6],afi_wdata[5],afi_wdata[4],afi_wdata[3],afi_wdata[2],afi_wdata[1],afi_wdata[0]}),
	.afiwdatavalid({afi_wdata_valid[4],afi_wdata_valid[3],afi_wdata_valid[2],afi_wdata_valid[1],afi_wdata_valid[0]}),
	.avladdress({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.avlwritedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfgaddlat({gnd,gnd,gnd,cfg_addlat[4],cfg_addlat[3],cfg_addlat[2],cfg_addlat[1],cfg_addlat[0]}),
	.cfgbankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth[2],cfg_bankaddrwidth[1],cfg_bankaddrwidth[0]}),
	.cfgcaswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat[3],cfg_caswrlat[2],cfg_caswrlat[1],cfg_caswrlat[0]}),
	.cfgcoladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth[4],cfg_coladdrwidth[3],cfg_coladdrwidth[2],cfg_coladdrwidth[1],cfg_coladdrwidth[0]}),
	.cfgcsaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth[2],cfg_csaddrwidth[1],cfg_csaddrwidth[0]}),
	.cfgdevicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth[3],cfg_devicewidth[2],cfg_devicewidth[1],cfg_devicewidth[0]}),
	.cfgdramconfig({gnd,gnd,gnd,cfg_dramconfig[20],cfg_dramconfig[19],cfg_dramconfig[18],cfg_dramconfig[17],cfg_dramconfig[16],cfg_dramconfig[15],cfg_dramconfig[14],cfg_dramconfig[13],cfg_dramconfig[12],cfg_dramconfig[11],cfg_dramconfig[10],cfg_dramconfig[9],cfg_dramconfig[8],cfg_dramconfig[7],cfg_dramconfig[6],cfg_dramconfig[5],cfg_dramconfig[4],
cfg_dramconfig[3],cfg_dramconfig[2],cfg_dramconfig[1],cfg_dramconfig[0]}),
	.cfginterfacewidth({cfg_interfacewidth[7],cfg_interfacewidth[6],cfg_interfacewidth[5],cfg_interfacewidth[4],cfg_interfacewidth[3],cfg_interfacewidth[2],cfg_interfacewidth[1],cfg_interfacewidth[0]}),
	.cfgrowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth[4],cfg_rowaddrwidth[3],cfg_rowaddrwidth[2],cfg_rowaddrwidth[1],cfg_rowaddrwidth[0]}),
	.cfgtcl({gnd,gnd,gnd,cfg_tcl[4],cfg_tcl[3],cfg_tcl[2],cfg_tcl[1],cfg_tcl[0]}),
	.cfgtmrd({gnd,gnd,gnd,gnd,cfg_tmrd[3],cfg_tmrd[2],cfg_tmrd[1],cfg_tmrd[0]}),
	.cfgtrefi({gnd,gnd,gnd,cfg_trefi[12],cfg_trefi[11],cfg_trefi[10],cfg_trefi[9],cfg_trefi[8],cfg_trefi[7],cfg_trefi[6],cfg_trefi[5],cfg_trefi[4],cfg_trefi[3],cfg_trefi[2],cfg_trefi[1],cfg_trefi[0]}),
	.cfgtrfc({cfg_trfc[7],cfg_trfc[6],cfg_trfc[5],cfg_trfc[4],cfg_trfc[3],cfg_trfc[2],cfg_trfc[1],cfg_trfc[0]}),
	.cfgtwr({gnd,gnd,gnd,gnd,cfg_twr[3],cfg_twr[2],cfg_twr[1],cfg_twr[0]}),
	.ddiophydqdin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] }),
	.ddiophydqslogicrdatavalid({vcc,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.iointaddraclr(16'b0000000000000000),
	.iointaddrdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointbaaclr(3'b000),
	.iointbadout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointcasndout({gnd,gnd,gnd,gnd}),
	.iointckdout({gnd,gnd,gnd,gnd}),
	.iointckeaclr(2'b00),
	.iointckedout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointckndout({gnd,gnd,gnd,gnd}),
	.iointcsnaclr(2'b00),
	.iointcsndout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdmdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iointdqsbdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsboe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicaclrfifoctrl(5'b00000),
	.iointdqslogicaclrpstamble(5'b00000),
	.iointdqslogicdqsena({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicfiforeset({gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincrdataen({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincwrptr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicoct({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicreadlatency({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointodtaclr(2'b00),
	.iointodtdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointrasndout({gnd,gnd,gnd,gnd}),
	.iointresetndout({gnd,gnd,gnd,gnd}),
	.iointwendout({gnd,gnd,gnd,gnd}),
	.aficalfail(afi_cal_fail),
	.aficalsuccess(afi_cal_success),
	.afirdatavalid(afi_rdata_valid[0]),
	.avlwaitrequest(),
	.ctlresetn(ctl_reset_n),
	.iointaficalfail(),
	.iointaficalsuccess(),
	.phyddiocasnaclr(),
	.phyddiorasnaclr(),
	.phyddioresetnaclr(),
	.phyddiowenaclr(),
	.phyresetn(),
	.afirdata(hphy_inst_AFIRDATA_bus),
	.afirlat(),
	.afiwlat(hphy_inst_AFIWLAT_bus),
	.avlreaddata(),
	.iointafirlat(),
	.iointafiwlat(),
	.iointdqdin(),
	.iointdqslogicrdatavalid(),
	.phyddioaddraclr(),
	.phyddioaddrdout(hphy_inst_PHYDDIOADDRDOUT_bus),
	.phyddiobaaclr(),
	.phyddiobadout(hphy_inst_PHYDDIOBADOUT_bus),
	.phyddiocasndout(hphy_inst_PHYDDIOCASNDOUT_bus),
	.phyddiockdout(hphy_inst_PHYDDIOCKDOUT_bus),
	.phyddiockeaclr(),
	.phyddiockedout(hphy_inst_PHYDDIOCKEDOUT_bus),
	.phyddiockndout(),
	.phyddiocsnaclr(),
	.phyddiocsndout(hphy_inst_PHYDDIOCSNDOUT_bus),
	.phyddiodmdout(hphy_inst_PHYDDIODMDOUT_bus),
	.phyddiodqdout(hphy_inst_PHYDDIODQDOUT_bus),
	.phyddiodqoe(hphy_inst_PHYDDIODQOE_bus),
	.phyddiodqsbdout(),
	.phyddiodqsboe(),
	.phyddiodqsdout(hphy_inst_PHYDDIODQSDOUT_bus),
	.phyddiodqslogicaclrfifoctrl(hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus),
	.phyddiodqslogicaclrpstamble(hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus),
	.phyddiodqslogicdqsena(hphy_inst_PHYDDIODQSLOGICDQSENA_bus),
	.phyddiodqslogicfiforeset(hphy_inst_PHYDDIODQSLOGICFIFORESET_bus),
	.phyddiodqslogicincrdataen(hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus),
	.phyddiodqslogicincwrptr(hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus),
	.phyddiodqslogicoct(hphy_inst_PHYDDIODQSLOGICOCT_bus),
	.phyddiodqslogicreadlatency(hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus),
	.phyddiodqsoe(hphy_inst_PHYDDIODQSOE_bus),
	.phyddioodtaclr(),
	.phyddioodtdout(hphy_inst_PHYDDIOODTDOUT_bus),
	.phyddiorasndout(hphy_inst_PHYDDIORASNDOUT_bus),
	.phyddioresetndout(hphy_inst_PHYDDIORESETNDOUT_bus),
	.phyddiowendout(hphy_inst_PHYDDIOWENDOUT_bus));
defparam hphy_inst.hphy_ac_ddr_disable = "true";
defparam hphy_inst.hphy_atpg_en = "false";
defparam hphy_inst.hphy_csr_pipelineglobalenable = "true";
defparam hphy_inst.hphy_datapath_ac_delay = "one_and_half_cycles";
defparam hphy_inst.hphy_datapath_delay = "one_cycle";
defparam hphy_inst.hphy_reset_delay_en = "false";
defparam hphy_inst.hphy_use_hphy = "true";
defparam hphy_inst.hphy_wrap_back_en = "false";
defparam hphy_inst.m_hphy_ac_rom_content = 1200'b100000011100000000000000000000100000011110000000000000000000010000000010000000010001110001010000000010000000010101110000010000000010010000000000000110010000000010100000001000011000010000000010110000000000000000010000001110000000010000000000010000000010000000010001101001010000000010000000010011101000010000000010100000000000000110010000000010010000001000011000010000000010110000000000000000110000011110000000000000000000111000011110000000000000000000110000011110000000000000000000010000011010000000000000000000010000011010110000000000000000010000001010000000010000000000010000010010000000000000000000011100100110000000000000000000011100100110110000000000000000011100100110000000000000001000011100100110110000000000001000111000111110000000000000000000111100111110000000000000000000111000011110000000000000000000011000000110000000000000000000011000100110000000000000000000010011010110000000000000000000010011010110110000000000000000010011010110000000000000001000010011010110110000000000001000110011011110000000000000000000010000010110000000000000001000010000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam hphy_inst.m_hphy_ac_rom_init_file = "hps_ac_rom.hex";
defparam hphy_inst.m_hphy_inst_rom_content = 2560'b1000000000000000000010000000011010000000000010000001100000000000100000100000000000001000001010000000000010000011000000000000100000111000000000001000000100000000000010000100100000000000100001010000000000001000010110000000000010000110000000000000100001000000000000000000100000000000000010000110100000000000000010001000000000001010011010000000100000000110100000000000000010010000000010000000011010000000000000001001100000000000101001101000000000001000011010000000100000000110100000000000000010110110100000001100110011101000000000001010111010000000100011001110100000000000101110001000000011101100100010000000000010100000100000001010110010001000100000000110100000000000110011100000000000001100110110000000000011100111000000000000000011000000000000100000110011100000001000001100111000000010000011001110000000100000110011100000000000001101000000000000000001101000000000000000011010000000000000000110100000000000000001101000000001100000111010000000011000010000100000000110000100001000000001100001000010000000000010100110100000000000100001101000000010000000011010000000000011001110000000000000110011011000000000001110011100000000000000001100000000000011000011001110000000110000110011100000001100001100111000000011000011001110000000000000110100000000000000000110100000000000000001101000000000000000011010000000000000000110100000000111000011101000000001110001000010000000011100010000100000000111000100001000000000001010011010000000000010000110100000001000000001101000000000000001000101011000000000000110110110001000000001101000000000000001000101101000000000000111111010000000000001111110100000001000011111101000010000001111111010000100000100001110100001000001000011101000010000010000111010000000000100010110100000000000011111101000000000000111111010000000101001111110100010000000011010000000010000001110100010000100000100001000100001000001000010001000010000010000100010000100000011110110100001000001000011101000010000010000111010000100000100001110100000001010011010000000010000001111111010000100000100001110100001000001000011101000010000010000111010000100000100000000100001000001000010001000010000010000100010000100000100001000100000000001000100000000000011000110100000000000100001101000000000001110011010000000100000000110100000000000000000000000000000001000000000000000000010100000000000000000110000000000000010000000000000000000000000000000100000000000100000001000000000001010000010000000000011000000100000001000000000001000000000001001000110000000000010000110100000000000101001101000000010000000011010000000010000001111000010001000000001101000000000000000000000000000;
defparam hphy_inst.m_hphy_inst_rom_init_file = "hps_inst_rom.hex";

endmodule

module system_hps_sdram_p0_acv_hard_io_pads (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	input_path_gen0read_fifo_out_01,
	input_path_gen0read_fifo_out_11,
	input_path_gen0read_fifo_out_21,
	input_path_gen0read_fifo_out_31,
	input_path_gen1read_fifo_out_01,
	input_path_gen1read_fifo_out_11,
	input_path_gen1read_fifo_out_21,
	input_path_gen1read_fifo_out_31,
	input_path_gen2read_fifo_out_01,
	input_path_gen2read_fifo_out_11,
	input_path_gen2read_fifo_out_21,
	input_path_gen2read_fifo_out_31,
	input_path_gen3read_fifo_out_01,
	input_path_gen3read_fifo_out_11,
	input_path_gen3read_fifo_out_21,
	input_path_gen3read_fifo_out_31,
	input_path_gen4read_fifo_out_01,
	input_path_gen4read_fifo_out_11,
	input_path_gen4read_fifo_out_21,
	input_path_gen4read_fifo_out_31,
	input_path_gen5read_fifo_out_01,
	input_path_gen5read_fifo_out_11,
	input_path_gen5read_fifo_out_21,
	input_path_gen5read_fifo_out_31,
	input_path_gen6read_fifo_out_01,
	input_path_gen6read_fifo_out_11,
	input_path_gen6read_fifo_out_21,
	input_path_gen6read_fifo_out_31,
	input_path_gen7read_fifo_out_01,
	input_path_gen7read_fifo_out_11,
	input_path_gen7read_fifo_out_21,
	input_path_gen7read_fifo_out_31,
	input_path_gen0read_fifo_out_02,
	input_path_gen0read_fifo_out_12,
	input_path_gen0read_fifo_out_22,
	input_path_gen0read_fifo_out_32,
	input_path_gen1read_fifo_out_02,
	input_path_gen1read_fifo_out_12,
	input_path_gen1read_fifo_out_22,
	input_path_gen1read_fifo_out_32,
	input_path_gen2read_fifo_out_02,
	input_path_gen2read_fifo_out_12,
	input_path_gen2read_fifo_out_22,
	input_path_gen2read_fifo_out_32,
	input_path_gen3read_fifo_out_02,
	input_path_gen3read_fifo_out_12,
	input_path_gen3read_fifo_out_22,
	input_path_gen3read_fifo_out_32,
	input_path_gen4read_fifo_out_02,
	input_path_gen4read_fifo_out_12,
	input_path_gen4read_fifo_out_22,
	input_path_gen4read_fifo_out_32,
	input_path_gen5read_fifo_out_02,
	input_path_gen5read_fifo_out_12,
	input_path_gen5read_fifo_out_22,
	input_path_gen5read_fifo_out_32,
	input_path_gen6read_fifo_out_02,
	input_path_gen6read_fifo_out_12,
	input_path_gen6read_fifo_out_22,
	input_path_gen6read_fifo_out_32,
	input_path_gen7read_fifo_out_02,
	input_path_gen7read_fifo_out_12,
	input_path_gen7read_fifo_out_22,
	input_path_gen7read_fifo_out_32,
	input_path_gen0read_fifo_out_03,
	input_path_gen0read_fifo_out_13,
	input_path_gen0read_fifo_out_23,
	input_path_gen0read_fifo_out_33,
	input_path_gen1read_fifo_out_03,
	input_path_gen1read_fifo_out_13,
	input_path_gen1read_fifo_out_23,
	input_path_gen1read_fifo_out_33,
	input_path_gen2read_fifo_out_03,
	input_path_gen2read_fifo_out_13,
	input_path_gen2read_fifo_out_23,
	input_path_gen2read_fifo_out_33,
	input_path_gen3read_fifo_out_03,
	input_path_gen3read_fifo_out_13,
	input_path_gen3read_fifo_out_23,
	input_path_gen3read_fifo_out_33,
	input_path_gen4read_fifo_out_03,
	input_path_gen4read_fifo_out_13,
	input_path_gen4read_fifo_out_23,
	input_path_gen4read_fifo_out_33,
	input_path_gen5read_fifo_out_03,
	input_path_gen5read_fifo_out_13,
	input_path_gen5read_fifo_out_23,
	input_path_gen5read_fifo_out_33,
	input_path_gen6read_fifo_out_03,
	input_path_gen6read_fifo_out_13,
	input_path_gen6read_fifo_out_23,
	input_path_gen6read_fifo_out_33,
	input_path_gen7read_fifo_out_03,
	input_path_gen7read_fifo_out_13,
	input_path_gen7read_fifo_out_23,
	input_path_gen7read_fifo_out_33,
	ddio_phy_dqslogic_rdatavalid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	input_path_gen0read_fifo_out_01;
output 	input_path_gen0read_fifo_out_11;
output 	input_path_gen0read_fifo_out_21;
output 	input_path_gen0read_fifo_out_31;
output 	input_path_gen1read_fifo_out_01;
output 	input_path_gen1read_fifo_out_11;
output 	input_path_gen1read_fifo_out_21;
output 	input_path_gen1read_fifo_out_31;
output 	input_path_gen2read_fifo_out_01;
output 	input_path_gen2read_fifo_out_11;
output 	input_path_gen2read_fifo_out_21;
output 	input_path_gen2read_fifo_out_31;
output 	input_path_gen3read_fifo_out_01;
output 	input_path_gen3read_fifo_out_11;
output 	input_path_gen3read_fifo_out_21;
output 	input_path_gen3read_fifo_out_31;
output 	input_path_gen4read_fifo_out_01;
output 	input_path_gen4read_fifo_out_11;
output 	input_path_gen4read_fifo_out_21;
output 	input_path_gen4read_fifo_out_31;
output 	input_path_gen5read_fifo_out_01;
output 	input_path_gen5read_fifo_out_11;
output 	input_path_gen5read_fifo_out_21;
output 	input_path_gen5read_fifo_out_31;
output 	input_path_gen6read_fifo_out_01;
output 	input_path_gen6read_fifo_out_11;
output 	input_path_gen6read_fifo_out_21;
output 	input_path_gen6read_fifo_out_31;
output 	input_path_gen7read_fifo_out_01;
output 	input_path_gen7read_fifo_out_11;
output 	input_path_gen7read_fifo_out_21;
output 	input_path_gen7read_fifo_out_31;
output 	input_path_gen0read_fifo_out_02;
output 	input_path_gen0read_fifo_out_12;
output 	input_path_gen0read_fifo_out_22;
output 	input_path_gen0read_fifo_out_32;
output 	input_path_gen1read_fifo_out_02;
output 	input_path_gen1read_fifo_out_12;
output 	input_path_gen1read_fifo_out_22;
output 	input_path_gen1read_fifo_out_32;
output 	input_path_gen2read_fifo_out_02;
output 	input_path_gen2read_fifo_out_12;
output 	input_path_gen2read_fifo_out_22;
output 	input_path_gen2read_fifo_out_32;
output 	input_path_gen3read_fifo_out_02;
output 	input_path_gen3read_fifo_out_12;
output 	input_path_gen3read_fifo_out_22;
output 	input_path_gen3read_fifo_out_32;
output 	input_path_gen4read_fifo_out_02;
output 	input_path_gen4read_fifo_out_12;
output 	input_path_gen4read_fifo_out_22;
output 	input_path_gen4read_fifo_out_32;
output 	input_path_gen5read_fifo_out_02;
output 	input_path_gen5read_fifo_out_12;
output 	input_path_gen5read_fifo_out_22;
output 	input_path_gen5read_fifo_out_32;
output 	input_path_gen6read_fifo_out_02;
output 	input_path_gen6read_fifo_out_12;
output 	input_path_gen6read_fifo_out_22;
output 	input_path_gen6read_fifo_out_32;
output 	input_path_gen7read_fifo_out_02;
output 	input_path_gen7read_fifo_out_12;
output 	input_path_gen7read_fifo_out_22;
output 	input_path_gen7read_fifo_out_32;
output 	input_path_gen0read_fifo_out_03;
output 	input_path_gen0read_fifo_out_13;
output 	input_path_gen0read_fifo_out_23;
output 	input_path_gen0read_fifo_out_33;
output 	input_path_gen1read_fifo_out_03;
output 	input_path_gen1read_fifo_out_13;
output 	input_path_gen1read_fifo_out_23;
output 	input_path_gen1read_fifo_out_33;
output 	input_path_gen2read_fifo_out_03;
output 	input_path_gen2read_fifo_out_13;
output 	input_path_gen2read_fifo_out_23;
output 	input_path_gen2read_fifo_out_33;
output 	input_path_gen3read_fifo_out_03;
output 	input_path_gen3read_fifo_out_13;
output 	input_path_gen3read_fifo_out_23;
output 	input_path_gen3read_fifo_out_33;
output 	input_path_gen4read_fifo_out_03;
output 	input_path_gen4read_fifo_out_13;
output 	input_path_gen4read_fifo_out_23;
output 	input_path_gen4read_fifo_out_33;
output 	input_path_gen5read_fifo_out_03;
output 	input_path_gen5read_fifo_out_13;
output 	input_path_gen5read_fifo_out_23;
output 	input_path_gen5read_fifo_out_33;
output 	input_path_gen6read_fifo_out_03;
output 	input_path_gen6read_fifo_out_13;
output 	input_path_gen6read_fifo_out_23;
output 	input_path_gen6read_fifo_out_33;
output 	input_path_gen7read_fifo_out_03;
output 	input_path_gen7read_fifo_out_13;
output 	input_path_gen7read_fifo_out_23;
output 	input_path_gen7read_fifo_out_33;
output 	[4:0] ddio_phy_dqslogic_rdatavalid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_hps_sdram_p0_altdqdqs_3 \dq_ddio[3].ubidir_dq_dqs (
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.phy_ddio_dmdout_12(phy_ddio_dmdout_12),
	.phy_ddio_dmdout_13(phy_ddio_dmdout_13),
	.phy_ddio_dmdout_14(phy_ddio_dmdout_14),
	.phy_ddio_dmdout_15(phy_ddio_dmdout_15),
	.phy_ddio_dqdout_108(phy_ddio_dqdout_108),
	.phy_ddio_dqdout_109(phy_ddio_dqdout_109),
	.phy_ddio_dqdout_110(phy_ddio_dqdout_110),
	.phy_ddio_dqdout_111(phy_ddio_dqdout_111),
	.phy_ddio_dqdout_112(phy_ddio_dqdout_112),
	.phy_ddio_dqdout_113(phy_ddio_dqdout_113),
	.phy_ddio_dqdout_114(phy_ddio_dqdout_114),
	.phy_ddio_dqdout_115(phy_ddio_dqdout_115),
	.phy_ddio_dqdout_116(phy_ddio_dqdout_116),
	.phy_ddio_dqdout_117(phy_ddio_dqdout_117),
	.phy_ddio_dqdout_118(phy_ddio_dqdout_118),
	.phy_ddio_dqdout_119(phy_ddio_dqdout_119),
	.phy_ddio_dqdout_120(phy_ddio_dqdout_120),
	.phy_ddio_dqdout_121(phy_ddio_dqdout_121),
	.phy_ddio_dqdout_122(phy_ddio_dqdout_122),
	.phy_ddio_dqdout_123(phy_ddio_dqdout_123),
	.phy_ddio_dqdout_124(phy_ddio_dqdout_124),
	.phy_ddio_dqdout_125(phy_ddio_dqdout_125),
	.phy_ddio_dqdout_126(phy_ddio_dqdout_126),
	.phy_ddio_dqdout_127(phy_ddio_dqdout_127),
	.phy_ddio_dqdout_128(phy_ddio_dqdout_128),
	.phy_ddio_dqdout_129(phy_ddio_dqdout_129),
	.phy_ddio_dqdout_130(phy_ddio_dqdout_130),
	.phy_ddio_dqdout_131(phy_ddio_dqdout_131),
	.phy_ddio_dqdout_132(phy_ddio_dqdout_132),
	.phy_ddio_dqdout_133(phy_ddio_dqdout_133),
	.phy_ddio_dqdout_134(phy_ddio_dqdout_134),
	.phy_ddio_dqdout_135(phy_ddio_dqdout_135),
	.phy_ddio_dqdout_136(phy_ddio_dqdout_136),
	.phy_ddio_dqdout_137(phy_ddio_dqdout_137),
	.phy_ddio_dqdout_138(phy_ddio_dqdout_138),
	.phy_ddio_dqdout_139(phy_ddio_dqdout_139),
	.phy_ddio_dqoe_54(phy_ddio_dqoe_54),
	.phy_ddio_dqoe_55(phy_ddio_dqoe_55),
	.phy_ddio_dqoe_56(phy_ddio_dqoe_56),
	.phy_ddio_dqoe_57(phy_ddio_dqoe_57),
	.phy_ddio_dqoe_58(phy_ddio_dqoe_58),
	.phy_ddio_dqoe_59(phy_ddio_dqoe_59),
	.phy_ddio_dqoe_60(phy_ddio_dqoe_60),
	.phy_ddio_dqoe_61(phy_ddio_dqoe_61),
	.phy_ddio_dqoe_62(phy_ddio_dqoe_62),
	.phy_ddio_dqoe_63(phy_ddio_dqoe_63),
	.phy_ddio_dqoe_64(phy_ddio_dqoe_64),
	.phy_ddio_dqoe_65(phy_ddio_dqoe_65),
	.phy_ddio_dqoe_66(phy_ddio_dqoe_66),
	.phy_ddio_dqoe_67(phy_ddio_dqoe_67),
	.phy_ddio_dqoe_68(phy_ddio_dqoe_68),
	.phy_ddio_dqoe_69(phy_ddio_dqoe_69),
	.phy_ddio_dqs_dout_12(phy_ddio_dqs_dout_12),
	.phy_ddio_dqs_dout_13(phy_ddio_dqs_dout_13),
	.phy_ddio_dqs_dout_14(phy_ddio_dqs_dout_14),
	.phy_ddio_dqs_dout_15(phy_ddio_dqs_dout_15),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.phy_ddio_dqslogic_aclr_pstamble_3(phy_ddio_dqslogic_aclr_pstamble_3),
	.phy_ddio_dqslogic_dqsena_6(phy_ddio_dqslogic_dqsena_6),
	.phy_ddio_dqslogic_dqsena_7(phy_ddio_dqslogic_dqsena_7),
	.phy_ddio_dqslogic_fiforeset_3(phy_ddio_dqslogic_fiforeset_3),
	.phy_ddio_dqslogic_incrdataen_6(phy_ddio_dqslogic_incrdataen_6),
	.phy_ddio_dqslogic_incrdataen_7(phy_ddio_dqslogic_incrdataen_7),
	.phy_ddio_dqslogic_incwrptr_6(phy_ddio_dqslogic_incwrptr_6),
	.phy_ddio_dqslogic_incwrptr_7(phy_ddio_dqslogic_incwrptr_7),
	.phy_ddio_dqslogic_oct_6(phy_ddio_dqslogic_oct_6),
	.phy_ddio_dqslogic_oct_7(phy_ddio_dqslogic_oct_7),
	.phy_ddio_dqslogic_readlatency_15(phy_ddio_dqslogic_readlatency_15),
	.phy_ddio_dqslogic_readlatency_16(phy_ddio_dqslogic_readlatency_16),
	.phy_ddio_dqslogic_readlatency_17(phy_ddio_dqslogic_readlatency_17),
	.phy_ddio_dqslogic_readlatency_18(phy_ddio_dqslogic_readlatency_18),
	.phy_ddio_dqslogic_readlatency_19(phy_ddio_dqslogic_readlatency_19),
	.phy_ddio_dqs_oe_6(phy_ddio_dqs_oe_6),
	.phy_ddio_dqs_oe_7(phy_ddio_dqs_oe_7),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_13),
	.delayed_oct(delayed_oct3),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_13),
	.os(os3),
	.os_bar(os_bar3),
	.diff_oe(diff_oe3),
	.diff_oe_bar(diff_oe_bar3),
	.diff_dtc(diff_dtc3),
	.diff_dtc_bar(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_03),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_13),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_23),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_33),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_03),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_13),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_23),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_33),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_03),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_13),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_23),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_33),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_03),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_13),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_23),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_33),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_03),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_13),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_23),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_33),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_03),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_13),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_23),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_33),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_03),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_13),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_23),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_33),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_03),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_13),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_23),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_33),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[3]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

system_hps_sdram_p0_altdqdqs_2 \dq_ddio[2].ubidir_dq_dqs (
	.dqsin(dqsin1),
	.pad_gen0raw_input(pad_gen0raw_input1),
	.pad_gen1raw_input(pad_gen1raw_input1),
	.pad_gen2raw_input(pad_gen2raw_input1),
	.pad_gen3raw_input(pad_gen3raw_input1),
	.pad_gen4raw_input(pad_gen4raw_input1),
	.pad_gen5raw_input(pad_gen5raw_input1),
	.pad_gen6raw_input(pad_gen6raw_input1),
	.pad_gen7raw_input(pad_gen7raw_input1),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out1),
	.phy_ddio_dmdout_8(phy_ddio_dmdout_8),
	.phy_ddio_dmdout_9(phy_ddio_dmdout_9),
	.phy_ddio_dmdout_10(phy_ddio_dmdout_10),
	.phy_ddio_dmdout_11(phy_ddio_dmdout_11),
	.phy_ddio_dqdout_72(phy_ddio_dqdout_72),
	.phy_ddio_dqdout_73(phy_ddio_dqdout_73),
	.phy_ddio_dqdout_74(phy_ddio_dqdout_74),
	.phy_ddio_dqdout_75(phy_ddio_dqdout_75),
	.phy_ddio_dqdout_76(phy_ddio_dqdout_76),
	.phy_ddio_dqdout_77(phy_ddio_dqdout_77),
	.phy_ddio_dqdout_78(phy_ddio_dqdout_78),
	.phy_ddio_dqdout_79(phy_ddio_dqdout_79),
	.phy_ddio_dqdout_80(phy_ddio_dqdout_80),
	.phy_ddio_dqdout_81(phy_ddio_dqdout_81),
	.phy_ddio_dqdout_82(phy_ddio_dqdout_82),
	.phy_ddio_dqdout_83(phy_ddio_dqdout_83),
	.phy_ddio_dqdout_84(phy_ddio_dqdout_84),
	.phy_ddio_dqdout_85(phy_ddio_dqdout_85),
	.phy_ddio_dqdout_86(phy_ddio_dqdout_86),
	.phy_ddio_dqdout_87(phy_ddio_dqdout_87),
	.phy_ddio_dqdout_88(phy_ddio_dqdout_88),
	.phy_ddio_dqdout_89(phy_ddio_dqdout_89),
	.phy_ddio_dqdout_90(phy_ddio_dqdout_90),
	.phy_ddio_dqdout_91(phy_ddio_dqdout_91),
	.phy_ddio_dqdout_92(phy_ddio_dqdout_92),
	.phy_ddio_dqdout_93(phy_ddio_dqdout_93),
	.phy_ddio_dqdout_94(phy_ddio_dqdout_94),
	.phy_ddio_dqdout_95(phy_ddio_dqdout_95),
	.phy_ddio_dqdout_96(phy_ddio_dqdout_96),
	.phy_ddio_dqdout_97(phy_ddio_dqdout_97),
	.phy_ddio_dqdout_98(phy_ddio_dqdout_98),
	.phy_ddio_dqdout_99(phy_ddio_dqdout_99),
	.phy_ddio_dqdout_100(phy_ddio_dqdout_100),
	.phy_ddio_dqdout_101(phy_ddio_dqdout_101),
	.phy_ddio_dqdout_102(phy_ddio_dqdout_102),
	.phy_ddio_dqdout_103(phy_ddio_dqdout_103),
	.phy_ddio_dqoe_36(phy_ddio_dqoe_36),
	.phy_ddio_dqoe_37(phy_ddio_dqoe_37),
	.phy_ddio_dqoe_38(phy_ddio_dqoe_38),
	.phy_ddio_dqoe_39(phy_ddio_dqoe_39),
	.phy_ddio_dqoe_40(phy_ddio_dqoe_40),
	.phy_ddio_dqoe_41(phy_ddio_dqoe_41),
	.phy_ddio_dqoe_42(phy_ddio_dqoe_42),
	.phy_ddio_dqoe_43(phy_ddio_dqoe_43),
	.phy_ddio_dqoe_44(phy_ddio_dqoe_44),
	.phy_ddio_dqoe_45(phy_ddio_dqoe_45),
	.phy_ddio_dqoe_46(phy_ddio_dqoe_46),
	.phy_ddio_dqoe_47(phy_ddio_dqoe_47),
	.phy_ddio_dqoe_48(phy_ddio_dqoe_48),
	.phy_ddio_dqoe_49(phy_ddio_dqoe_49),
	.phy_ddio_dqoe_50(phy_ddio_dqoe_50),
	.phy_ddio_dqoe_51(phy_ddio_dqoe_51),
	.phy_ddio_dqs_dout_8(phy_ddio_dqs_dout_8),
	.phy_ddio_dqs_dout_9(phy_ddio_dqs_dout_9),
	.phy_ddio_dqs_dout_10(phy_ddio_dqs_dout_10),
	.phy_ddio_dqs_dout_11(phy_ddio_dqs_dout_11),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.phy_ddio_dqslogic_aclr_pstamble_2(phy_ddio_dqslogic_aclr_pstamble_2),
	.phy_ddio_dqslogic_dqsena_4(phy_ddio_dqslogic_dqsena_4),
	.phy_ddio_dqslogic_dqsena_5(phy_ddio_dqslogic_dqsena_5),
	.phy_ddio_dqslogic_fiforeset_2(phy_ddio_dqslogic_fiforeset_2),
	.phy_ddio_dqslogic_incrdataen_4(phy_ddio_dqslogic_incrdataen_4),
	.phy_ddio_dqslogic_incrdataen_5(phy_ddio_dqslogic_incrdataen_5),
	.phy_ddio_dqslogic_incwrptr_4(phy_ddio_dqslogic_incwrptr_4),
	.phy_ddio_dqslogic_incwrptr_5(phy_ddio_dqslogic_incwrptr_5),
	.phy_ddio_dqslogic_oct_4(phy_ddio_dqslogic_oct_4),
	.phy_ddio_dqslogic_oct_5(phy_ddio_dqslogic_oct_5),
	.phy_ddio_dqslogic_readlatency_10(phy_ddio_dqslogic_readlatency_10),
	.phy_ddio_dqslogic_readlatency_11(phy_ddio_dqslogic_readlatency_11),
	.phy_ddio_dqslogic_readlatency_12(phy_ddio_dqslogic_readlatency_12),
	.phy_ddio_dqslogic_readlatency_13(phy_ddio_dqslogic_readlatency_13),
	.phy_ddio_dqslogic_readlatency_14(phy_ddio_dqslogic_readlatency_14),
	.phy_ddio_dqs_oe_4(phy_ddio_dqs_oe_4),
	.phy_ddio_dqs_oe_5(phy_ddio_dqs_oe_5),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_12),
	.delayed_oct(delayed_oct2),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_12),
	.os(os2),
	.os_bar(os_bar2),
	.diff_oe(diff_oe2),
	.diff_oe_bar(diff_oe_bar2),
	.diff_dtc(diff_dtc2),
	.diff_dtc_bar(diff_dtc_bar2),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_02),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_12),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_22),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_32),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_02),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_12),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_22),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_32),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_02),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_12),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_22),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_32),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_02),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_12),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_22),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_32),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_02),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_12),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_22),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_32),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_02),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_12),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_22),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_32),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_02),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_12),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_22),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_32),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_02),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_12),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_22),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_32),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[2]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

system_hps_sdram_p0_altdqdqs_1 \dq_ddio[1].ubidir_dq_dqs (
	.dqsin(dqsin2),
	.pad_gen0raw_input(pad_gen0raw_input2),
	.pad_gen1raw_input(pad_gen1raw_input2),
	.pad_gen2raw_input(pad_gen2raw_input2),
	.pad_gen3raw_input(pad_gen3raw_input2),
	.pad_gen4raw_input(pad_gen4raw_input2),
	.pad_gen5raw_input(pad_gen5raw_input2),
	.pad_gen6raw_input(pad_gen6raw_input2),
	.pad_gen7raw_input(pad_gen7raw_input2),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out2),
	.phy_ddio_dmdout_4(phy_ddio_dmdout_4),
	.phy_ddio_dmdout_5(phy_ddio_dmdout_5),
	.phy_ddio_dmdout_6(phy_ddio_dmdout_6),
	.phy_ddio_dmdout_7(phy_ddio_dmdout_7),
	.phy_ddio_dqdout_36(phy_ddio_dqdout_36),
	.phy_ddio_dqdout_37(phy_ddio_dqdout_37),
	.phy_ddio_dqdout_38(phy_ddio_dqdout_38),
	.phy_ddio_dqdout_39(phy_ddio_dqdout_39),
	.phy_ddio_dqdout_40(phy_ddio_dqdout_40),
	.phy_ddio_dqdout_41(phy_ddio_dqdout_41),
	.phy_ddio_dqdout_42(phy_ddio_dqdout_42),
	.phy_ddio_dqdout_43(phy_ddio_dqdout_43),
	.phy_ddio_dqdout_44(phy_ddio_dqdout_44),
	.phy_ddio_dqdout_45(phy_ddio_dqdout_45),
	.phy_ddio_dqdout_46(phy_ddio_dqdout_46),
	.phy_ddio_dqdout_47(phy_ddio_dqdout_47),
	.phy_ddio_dqdout_48(phy_ddio_dqdout_48),
	.phy_ddio_dqdout_49(phy_ddio_dqdout_49),
	.phy_ddio_dqdout_50(phy_ddio_dqdout_50),
	.phy_ddio_dqdout_51(phy_ddio_dqdout_51),
	.phy_ddio_dqdout_52(phy_ddio_dqdout_52),
	.phy_ddio_dqdout_53(phy_ddio_dqdout_53),
	.phy_ddio_dqdout_54(phy_ddio_dqdout_54),
	.phy_ddio_dqdout_55(phy_ddio_dqdout_55),
	.phy_ddio_dqdout_56(phy_ddio_dqdout_56),
	.phy_ddio_dqdout_57(phy_ddio_dqdout_57),
	.phy_ddio_dqdout_58(phy_ddio_dqdout_58),
	.phy_ddio_dqdout_59(phy_ddio_dqdout_59),
	.phy_ddio_dqdout_60(phy_ddio_dqdout_60),
	.phy_ddio_dqdout_61(phy_ddio_dqdout_61),
	.phy_ddio_dqdout_62(phy_ddio_dqdout_62),
	.phy_ddio_dqdout_63(phy_ddio_dqdout_63),
	.phy_ddio_dqdout_64(phy_ddio_dqdout_64),
	.phy_ddio_dqdout_65(phy_ddio_dqdout_65),
	.phy_ddio_dqdout_66(phy_ddio_dqdout_66),
	.phy_ddio_dqdout_67(phy_ddio_dqdout_67),
	.phy_ddio_dqoe_18(phy_ddio_dqoe_18),
	.phy_ddio_dqoe_19(phy_ddio_dqoe_19),
	.phy_ddio_dqoe_20(phy_ddio_dqoe_20),
	.phy_ddio_dqoe_21(phy_ddio_dqoe_21),
	.phy_ddio_dqoe_22(phy_ddio_dqoe_22),
	.phy_ddio_dqoe_23(phy_ddio_dqoe_23),
	.phy_ddio_dqoe_24(phy_ddio_dqoe_24),
	.phy_ddio_dqoe_25(phy_ddio_dqoe_25),
	.phy_ddio_dqoe_26(phy_ddio_dqoe_26),
	.phy_ddio_dqoe_27(phy_ddio_dqoe_27),
	.phy_ddio_dqoe_28(phy_ddio_dqoe_28),
	.phy_ddio_dqoe_29(phy_ddio_dqoe_29),
	.phy_ddio_dqoe_30(phy_ddio_dqoe_30),
	.phy_ddio_dqoe_31(phy_ddio_dqoe_31),
	.phy_ddio_dqoe_32(phy_ddio_dqoe_32),
	.phy_ddio_dqoe_33(phy_ddio_dqoe_33),
	.phy_ddio_dqs_dout_4(phy_ddio_dqs_dout_4),
	.phy_ddio_dqs_dout_5(phy_ddio_dqs_dout_5),
	.phy_ddio_dqs_dout_6(phy_ddio_dqs_dout_6),
	.phy_ddio_dqs_dout_7(phy_ddio_dqs_dout_7),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.phy_ddio_dqslogic_aclr_pstamble_1(phy_ddio_dqslogic_aclr_pstamble_1),
	.phy_ddio_dqslogic_dqsena_2(phy_ddio_dqslogic_dqsena_2),
	.phy_ddio_dqslogic_dqsena_3(phy_ddio_dqslogic_dqsena_3),
	.phy_ddio_dqslogic_fiforeset_1(phy_ddio_dqslogic_fiforeset_1),
	.phy_ddio_dqslogic_incrdataen_2(phy_ddio_dqslogic_incrdataen_2),
	.phy_ddio_dqslogic_incrdataen_3(phy_ddio_dqslogic_incrdataen_3),
	.phy_ddio_dqslogic_incwrptr_2(phy_ddio_dqslogic_incwrptr_2),
	.phy_ddio_dqslogic_incwrptr_3(phy_ddio_dqslogic_incwrptr_3),
	.phy_ddio_dqslogic_oct_2(phy_ddio_dqslogic_oct_2),
	.phy_ddio_dqslogic_oct_3(phy_ddio_dqslogic_oct_3),
	.phy_ddio_dqslogic_readlatency_5(phy_ddio_dqslogic_readlatency_5),
	.phy_ddio_dqslogic_readlatency_6(phy_ddio_dqslogic_readlatency_6),
	.phy_ddio_dqslogic_readlatency_7(phy_ddio_dqslogic_readlatency_7),
	.phy_ddio_dqslogic_readlatency_8(phy_ddio_dqslogic_readlatency_8),
	.phy_ddio_dqslogic_readlatency_9(phy_ddio_dqslogic_readlatency_9),
	.phy_ddio_dqs_oe_2(phy_ddio_dqs_oe_2),
	.phy_ddio_dqs_oe_3(phy_ddio_dqs_oe_3),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_11),
	.delayed_oct(delayed_oct1),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_11),
	.os(os1),
	.os_bar(os_bar1),
	.diff_oe(diff_oe1),
	.diff_oe_bar(diff_oe_bar1),
	.diff_dtc(diff_dtc1),
	.diff_dtc_bar(diff_dtc_bar1),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_01),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_11),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_21),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_31),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_01),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_11),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_21),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_31),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_01),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_11),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_21),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_31),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_01),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_11),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_21),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_31),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_01),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_11),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_21),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_31),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_01),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_11),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_21),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_31),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_01),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_11),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_21),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_31),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_01),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_11),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_21),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_31),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[1]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

system_hps_sdram_p0_altdqdqs \dq_ddio[0].ubidir_dq_dqs (
	.dqsin(dqsin3),
	.pad_gen0raw_input(pad_gen0raw_input3),
	.pad_gen1raw_input(pad_gen1raw_input3),
	.pad_gen2raw_input(pad_gen2raw_input3),
	.pad_gen3raw_input(pad_gen3raw_input3),
	.pad_gen4raw_input(pad_gen4raw_input3),
	.pad_gen5raw_input(pad_gen5raw_input3),
	.pad_gen6raw_input(pad_gen6raw_input3),
	.pad_gen7raw_input(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out3),
	.phy_ddio_dmdout_0(phy_ddio_dmdout_0),
	.phy_ddio_dmdout_1(phy_ddio_dmdout_1),
	.phy_ddio_dmdout_2(phy_ddio_dmdout_2),
	.phy_ddio_dmdout_3(phy_ddio_dmdout_3),
	.phy_ddio_dqdout_0(phy_ddio_dqdout_0),
	.phy_ddio_dqdout_1(phy_ddio_dqdout_1),
	.phy_ddio_dqdout_2(phy_ddio_dqdout_2),
	.phy_ddio_dqdout_3(phy_ddio_dqdout_3),
	.phy_ddio_dqdout_4(phy_ddio_dqdout_4),
	.phy_ddio_dqdout_5(phy_ddio_dqdout_5),
	.phy_ddio_dqdout_6(phy_ddio_dqdout_6),
	.phy_ddio_dqdout_7(phy_ddio_dqdout_7),
	.phy_ddio_dqdout_8(phy_ddio_dqdout_8),
	.phy_ddio_dqdout_9(phy_ddio_dqdout_9),
	.phy_ddio_dqdout_10(phy_ddio_dqdout_10),
	.phy_ddio_dqdout_11(phy_ddio_dqdout_11),
	.phy_ddio_dqdout_12(phy_ddio_dqdout_12),
	.phy_ddio_dqdout_13(phy_ddio_dqdout_13),
	.phy_ddio_dqdout_14(phy_ddio_dqdout_14),
	.phy_ddio_dqdout_15(phy_ddio_dqdout_15),
	.phy_ddio_dqdout_16(phy_ddio_dqdout_16),
	.phy_ddio_dqdout_17(phy_ddio_dqdout_17),
	.phy_ddio_dqdout_18(phy_ddio_dqdout_18),
	.phy_ddio_dqdout_19(phy_ddio_dqdout_19),
	.phy_ddio_dqdout_20(phy_ddio_dqdout_20),
	.phy_ddio_dqdout_21(phy_ddio_dqdout_21),
	.phy_ddio_dqdout_22(phy_ddio_dqdout_22),
	.phy_ddio_dqdout_23(phy_ddio_dqdout_23),
	.phy_ddio_dqdout_24(phy_ddio_dqdout_24),
	.phy_ddio_dqdout_25(phy_ddio_dqdout_25),
	.phy_ddio_dqdout_26(phy_ddio_dqdout_26),
	.phy_ddio_dqdout_27(phy_ddio_dqdout_27),
	.phy_ddio_dqdout_28(phy_ddio_dqdout_28),
	.phy_ddio_dqdout_29(phy_ddio_dqdout_29),
	.phy_ddio_dqdout_30(phy_ddio_dqdout_30),
	.phy_ddio_dqdout_31(phy_ddio_dqdout_31),
	.phy_ddio_dqoe_0(phy_ddio_dqoe_0),
	.phy_ddio_dqoe_1(phy_ddio_dqoe_1),
	.phy_ddio_dqoe_2(phy_ddio_dqoe_2),
	.phy_ddio_dqoe_3(phy_ddio_dqoe_3),
	.phy_ddio_dqoe_4(phy_ddio_dqoe_4),
	.phy_ddio_dqoe_5(phy_ddio_dqoe_5),
	.phy_ddio_dqoe_6(phy_ddio_dqoe_6),
	.phy_ddio_dqoe_7(phy_ddio_dqoe_7),
	.phy_ddio_dqoe_8(phy_ddio_dqoe_8),
	.phy_ddio_dqoe_9(phy_ddio_dqoe_9),
	.phy_ddio_dqoe_10(phy_ddio_dqoe_10),
	.phy_ddio_dqoe_11(phy_ddio_dqoe_11),
	.phy_ddio_dqoe_12(phy_ddio_dqoe_12),
	.phy_ddio_dqoe_13(phy_ddio_dqoe_13),
	.phy_ddio_dqoe_14(phy_ddio_dqoe_14),
	.phy_ddio_dqoe_15(phy_ddio_dqoe_15),
	.phy_ddio_dqs_dout_0(phy_ddio_dqs_dout_0),
	.phy_ddio_dqs_dout_1(phy_ddio_dqs_dout_1),
	.phy_ddio_dqs_dout_2(phy_ddio_dqs_dout_2),
	.phy_ddio_dqs_dout_3(phy_ddio_dqs_dout_3),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.phy_ddio_dqslogic_aclr_pstamble_0(phy_ddio_dqslogic_aclr_pstamble_0),
	.phy_ddio_dqslogic_dqsena_0(phy_ddio_dqslogic_dqsena_0),
	.phy_ddio_dqslogic_dqsena_1(phy_ddio_dqslogic_dqsena_1),
	.phy_ddio_dqslogic_fiforeset_0(phy_ddio_dqslogic_fiforeset_0),
	.phy_ddio_dqslogic_incrdataen_0(phy_ddio_dqslogic_incrdataen_0),
	.phy_ddio_dqslogic_incrdataen_1(phy_ddio_dqslogic_incrdataen_1),
	.phy_ddio_dqslogic_incwrptr_0(phy_ddio_dqslogic_incwrptr_0),
	.phy_ddio_dqslogic_incwrptr_1(phy_ddio_dqslogic_incwrptr_1),
	.phy_ddio_dqslogic_oct_0(phy_ddio_dqslogic_oct_0),
	.phy_ddio_dqslogic_oct_1(phy_ddio_dqslogic_oct_1),
	.phy_ddio_dqslogic_readlatency_0(phy_ddio_dqslogic_readlatency_0),
	.phy_ddio_dqslogic_readlatency_1(phy_ddio_dqslogic_readlatency_1),
	.phy_ddio_dqslogic_readlatency_2(phy_ddio_dqslogic_readlatency_2),
	.phy_ddio_dqslogic_readlatency_3(phy_ddio_dqslogic_readlatency_3),
	.phy_ddio_dqslogic_readlatency_4(phy_ddio_dqslogic_readlatency_4),
	.phy_ddio_dqs_oe_0(phy_ddio_dqs_oe_0),
	.phy_ddio_dqs_oe_1(phy_ddio_dqs_oe_1),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_0),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_1),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_2),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_3),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_0),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_1),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_2),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_3),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_0),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_1),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_2),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_3),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_0),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_1),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_2),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_3),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_0),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_1),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_2),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_3),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_0),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_1),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_2),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_3),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_0),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_1),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_2),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_3),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_0),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_1),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_2),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_3),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[0]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

system_hps_sdram_p0_acv_hard_addr_cmd_pads uaddr_cmd_pads(
	.afi_clk(afi_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(phy_ddio_address_0),
	.phy_ddio_address_1(phy_ddio_address_1),
	.phy_ddio_address_2(phy_ddio_address_2),
	.phy_ddio_address_3(phy_ddio_address_3),
	.phy_ddio_address_4(phy_ddio_address_4),
	.phy_ddio_address_5(phy_ddio_address_5),
	.phy_ddio_address_6(phy_ddio_address_6),
	.phy_ddio_address_7(phy_ddio_address_7),
	.phy_ddio_address_8(phy_ddio_address_8),
	.phy_ddio_address_9(phy_ddio_address_9),
	.phy_ddio_address_10(phy_ddio_address_10),
	.phy_ddio_address_11(phy_ddio_address_11),
	.phy_ddio_address_12(phy_ddio_address_12),
	.phy_ddio_address_13(phy_ddio_address_13),
	.phy_ddio_address_14(phy_ddio_address_14),
	.phy_ddio_address_15(phy_ddio_address_15),
	.phy_ddio_address_16(phy_ddio_address_16),
	.phy_ddio_address_17(phy_ddio_address_17),
	.phy_ddio_address_18(phy_ddio_address_18),
	.phy_ddio_address_19(phy_ddio_address_19),
	.phy_ddio_address_20(phy_ddio_address_20),
	.phy_ddio_address_21(phy_ddio_address_21),
	.phy_ddio_address_22(phy_ddio_address_22),
	.phy_ddio_address_23(phy_ddio_address_23),
	.phy_ddio_address_24(phy_ddio_address_24),
	.phy_ddio_address_25(phy_ddio_address_25),
	.phy_ddio_address_26(phy_ddio_address_26),
	.phy_ddio_address_27(phy_ddio_address_27),
	.phy_ddio_address_28(phy_ddio_address_28),
	.phy_ddio_address_29(phy_ddio_address_29),
	.phy_ddio_address_30(phy_ddio_address_30),
	.phy_ddio_address_31(phy_ddio_address_31),
	.phy_ddio_address_32(phy_ddio_address_32),
	.phy_ddio_address_33(phy_ddio_address_33),
	.phy_ddio_address_34(phy_ddio_address_34),
	.phy_ddio_address_35(phy_ddio_address_35),
	.phy_ddio_address_36(phy_ddio_address_36),
	.phy_ddio_address_37(phy_ddio_address_37),
	.phy_ddio_address_38(phy_ddio_address_38),
	.phy_ddio_address_39(phy_ddio_address_39),
	.phy_ddio_address_40(phy_ddio_address_40),
	.phy_ddio_address_41(phy_ddio_address_41),
	.phy_ddio_address_42(phy_ddio_address_42),
	.phy_ddio_address_43(phy_ddio_address_43),
	.phy_ddio_address_44(phy_ddio_address_44),
	.phy_ddio_address_45(phy_ddio_address_45),
	.phy_ddio_address_46(phy_ddio_address_46),
	.phy_ddio_address_47(phy_ddio_address_47),
	.phy_ddio_address_48(phy_ddio_address_48),
	.phy_ddio_address_49(phy_ddio_address_49),
	.phy_ddio_address_50(phy_ddio_address_50),
	.phy_ddio_address_51(phy_ddio_address_51),
	.phy_ddio_address_52(phy_ddio_address_52),
	.phy_ddio_address_53(phy_ddio_address_53),
	.phy_ddio_address_54(phy_ddio_address_54),
	.phy_ddio_address_55(phy_ddio_address_55),
	.phy_ddio_address_56(phy_ddio_address_56),
	.phy_ddio_address_57(phy_ddio_address_57),
	.phy_ddio_address_58(phy_ddio_address_58),
	.phy_ddio_address_59(phy_ddio_address_59),
	.phy_ddio_bank_0(phy_ddio_bank_0),
	.phy_ddio_bank_1(phy_ddio_bank_1),
	.phy_ddio_bank_2(phy_ddio_bank_2),
	.phy_ddio_bank_3(phy_ddio_bank_3),
	.phy_ddio_bank_4(phy_ddio_bank_4),
	.phy_ddio_bank_5(phy_ddio_bank_5),
	.phy_ddio_bank_6(phy_ddio_bank_6),
	.phy_ddio_bank_7(phy_ddio_bank_7),
	.phy_ddio_bank_8(phy_ddio_bank_8),
	.phy_ddio_bank_9(phy_ddio_bank_9),
	.phy_ddio_bank_10(phy_ddio_bank_10),
	.phy_ddio_bank_11(phy_ddio_bank_11),
	.phy_ddio_cas_n_0(phy_ddio_cas_n_0),
	.phy_ddio_cas_n_1(phy_ddio_cas_n_1),
	.phy_ddio_cas_n_2(phy_ddio_cas_n_2),
	.phy_ddio_cas_n_3(phy_ddio_cas_n_3),
	.phy_ddio_ck_0(phy_ddio_ck_0),
	.phy_ddio_ck_1(phy_ddio_ck_1),
	.phy_ddio_cke_0(phy_ddio_cke_0),
	.phy_ddio_cke_1(phy_ddio_cke_1),
	.phy_ddio_cke_2(phy_ddio_cke_2),
	.phy_ddio_cke_3(phy_ddio_cke_3),
	.phy_ddio_cs_n_0(phy_ddio_cs_n_0),
	.phy_ddio_cs_n_1(phy_ddio_cs_n_1),
	.phy_ddio_cs_n_2(phy_ddio_cs_n_2),
	.phy_ddio_cs_n_3(phy_ddio_cs_n_3),
	.phy_ddio_odt_0(phy_ddio_odt_0),
	.phy_ddio_odt_1(phy_ddio_odt_1),
	.phy_ddio_odt_2(phy_ddio_odt_2),
	.phy_ddio_odt_3(phy_ddio_odt_3),
	.phy_ddio_ras_n_0(phy_ddio_ras_n_0),
	.phy_ddio_ras_n_1(phy_ddio_ras_n_1),
	.phy_ddio_ras_n_2(phy_ddio_ras_n_2),
	.phy_ddio_ras_n_3(phy_ddio_ras_n_3),
	.phy_ddio_reset_n_0(phy_ddio_reset_n_0),
	.phy_ddio_reset_n_1(phy_ddio_reset_n_1),
	.phy_ddio_reset_n_2(phy_ddio_reset_n_2),
	.phy_ddio_reset_n_3(phy_ddio_reset_n_3),
	.phy_ddio_we_n_0(phy_ddio_we_n_0),
	.phy_ddio_we_n_1(phy_ddio_we_n_1),
	.phy_ddio_we_n_2(phy_ddio_we_n_2),
	.phy_ddio_we_n_3(phy_ddio_we_n_3),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6));

endmodule

module system_hps_sdram_p0_acv_hard_addr_cmd_pads (
	afi_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6)/* synthesis synthesis_greybox=0 */;
input 	afi_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_gen[0].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[1].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[2].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[3].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[4].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[5].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[6].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[7].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[8].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[9].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[10].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[11].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[12].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[13].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[14].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[15].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[16].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[17].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[19].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[18].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[21].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[22].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[23].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[24].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[20].acv_ac_ldc|adc_clk_cps ;
wire \clock_gen[0].umem_ck_pad|auto_generated|dataout[0] ;
wire \mem_ck_source[0] ;
wire \clock_gen[0].leveled_dqs_clocks[0] ;
wire \clock_gen[0].leveled_dqs_clocks[1] ;
wire \clock_gen[0].leveled_dqs_clocks[2] ;
wire \clock_gen[0].leveled_dqs_clocks[3] ;

wire [3:0] \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ;

assign \clock_gen[0].leveled_dqs_clocks[0]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [0];
assign \clock_gen[0].leveled_dqs_clocks[1]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [1];
assign \clock_gen[0].leveled_dqs_clocks[2]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [2];
assign \clock_gen[0].leveled_dqs_clocks[3]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [3];

system_hps_sdram_p0_clock_pair_generator \clock_gen[0].uclk_generator (
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.datain({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }));

system_altddio_out_1 \clock_gen[0].umem_ck_pad (
	.dataout({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }),
	.datain_h({phy_ddio_ck_0}),
	.datain_l({phy_ddio_ck_1}),
	.outclock(\mem_ck_source[0] ));

system_hps_sdram_p0_generic_ddio_3 ureset_n_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk}),
	.dataout({dataout_unconnected_wire_14,dataout_unconnected_wire_13,dataout_unconnected_wire_12,dataout_unconnected_wire_11,dataout_unconnected_wire_10,dataout_unconnected_wire_9,dataout_unconnected_wire_8,dataout_unconnected_wire_7,dataout_unconnected_wire_6,
dataout_unconnected_wire_5,dataout_unconnected_wire_4,dataout_unconnected_wire_3,dataout_unconnected_wire_2,dataout_unconnected_wire_1,dataout_03}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[24].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_reset_n_3,phy_ddio_reset_n_2,phy_ddio_reset_n_1,phy_ddio_reset_n_0}));

system_hps_sdram_p0_generic_ddio_2 ucmd_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_1,dataout_unconnected_wire_13_1,dataout_unconnected_wire_12_1,dataout_unconnected_wire_11_1,dataout_unconnected_wire_10_1,dataout_unconnected_wire_9_1,dataout_unconnected_wire_8_1,dataout_unconnected_wire_7_1,
dataout_unconnected_wire_6_1,dataout_51,dataout_41,dataout_31,dataout_22,dataout_16,dataout_02}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[23].acv_ac_ldc|adc_clk_cps ,\address_gen[22].acv_ac_ldc|adc_clk_cps ,\address_gen[21].acv_ac_ldc|adc_clk_cps ,\address_gen[20].acv_ac_ldc|adc_clk_cps ,\address_gen[19].acv_ac_ldc|adc_clk_cps ,
\address_gen[18].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_we_n_3,phy_ddio_we_n_2,phy_ddio_we_n_1,phy_ddio_we_n_0,phy_ddio_cas_n_3,phy_ddio_cas_n_2,phy_ddio_cas_n_1,phy_ddio_cas_n_0,phy_ddio_ras_n_3,
phy_ddio_ras_n_2,phy_ddio_ras_n_1,phy_ddio_ras_n_0,phy_ddio_odt_3,phy_ddio_odt_2,phy_ddio_odt_1,phy_ddio_odt_0,phy_ddio_cke_3,phy_ddio_cke_2,phy_ddio_cke_1,phy_ddio_cke_0,phy_ddio_cs_n_3,phy_ddio_cs_n_2,phy_ddio_cs_n_1,phy_ddio_cs_n_0}));

system_hps_sdram_p0_generic_ddio_1 ubank_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_2,dataout_unconnected_wire_13_2,dataout_unconnected_wire_12_2,dataout_unconnected_wire_11_2,dataout_unconnected_wire_10_2,dataout_unconnected_wire_9_2,dataout_unconnected_wire_8_2,dataout_unconnected_wire_7_2,
dataout_unconnected_wire_6_2,dataout_unconnected_wire_5_1,dataout_unconnected_wire_4_1,dataout_unconnected_wire_3_1,dataout_21,dataout_15,dataout_01}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[17].acv_ac_ldc|adc_clk_cps ,\address_gen[16].acv_ac_ldc|adc_clk_cps ,\address_gen[15].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_bank_11,phy_ddio_bank_10,phy_ddio_bank_9,phy_ddio_bank_8,phy_ddio_bank_7,phy_ddio_bank_6,phy_ddio_bank_5,
phy_ddio_bank_4,phy_ddio_bank_3,phy_ddio_bank_2,phy_ddio_bank_1,phy_ddio_bank_0}));

system_hps_sdram_p0_generic_ddio uaddress_pad(
	.clk_hr({afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_14,dataout_13,dataout_12,dataout_11,dataout_10,dataout_9,dataout_8,dataout_7,dataout_6,dataout_5,dataout_4,dataout_3,dataout_2,dataout_1,dataout_0}),
	.clk_fr({\address_gen[14].acv_ac_ldc|adc_clk_cps ,\address_gen[13].acv_ac_ldc|adc_clk_cps ,\address_gen[12].acv_ac_ldc|adc_clk_cps ,\address_gen[11].acv_ac_ldc|adc_clk_cps ,\address_gen[10].acv_ac_ldc|adc_clk_cps ,\address_gen[9].acv_ac_ldc|adc_clk_cps ,
\address_gen[8].acv_ac_ldc|adc_clk_cps ,\address_gen[7].acv_ac_ldc|adc_clk_cps ,\address_gen[6].acv_ac_ldc|adc_clk_cps ,\address_gen[5].acv_ac_ldc|adc_clk_cps ,\address_gen[4].acv_ac_ldc|adc_clk_cps ,\address_gen[3].acv_ac_ldc|adc_clk_cps ,
\address_gen[2].acv_ac_ldc|adc_clk_cps ,\address_gen[1].acv_ac_ldc|adc_clk_cps ,\address_gen[0].acv_ac_ldc|adc_clk_cps }),
	.datain({phy_ddio_address_59,phy_ddio_address_58,phy_ddio_address_57,phy_ddio_address_56,phy_ddio_address_55,phy_ddio_address_54,phy_ddio_address_53,phy_ddio_address_52,phy_ddio_address_51,phy_ddio_address_50,phy_ddio_address_49,phy_ddio_address_48,phy_ddio_address_47,
phy_ddio_address_46,phy_ddio_address_45,phy_ddio_address_44,phy_ddio_address_43,phy_ddio_address_42,phy_ddio_address_41,phy_ddio_address_40,phy_ddio_address_39,phy_ddio_address_38,phy_ddio_address_37,phy_ddio_address_36,phy_ddio_address_35,phy_ddio_address_34,
phy_ddio_address_33,phy_ddio_address_32,phy_ddio_address_31,phy_ddio_address_30,phy_ddio_address_29,phy_ddio_address_28,phy_ddio_address_27,phy_ddio_address_26,phy_ddio_address_25,phy_ddio_address_24,phy_ddio_address_23,phy_ddio_address_22,phy_ddio_address_21,
phy_ddio_address_20,phy_ddio_address_19,phy_ddio_address_18,phy_ddio_address_17,phy_ddio_address_16,phy_ddio_address_15,phy_ddio_address_14,phy_ddio_address_13,phy_ddio_address_12,phy_ddio_address_11,phy_ddio_address_10,phy_ddio_address_9,phy_ddio_address_8,
phy_ddio_address_7,phy_ddio_address_6,phy_ddio_address_5,phy_ddio_address_4,phy_ddio_address_3,phy_ddio_address_2,phy_ddio_address_1,phy_ddio_address_0}));

system_hps_sdram_p0_acv_ldc_16 \address_gen[24].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[24].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_15 \address_gen[23].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[23].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_14 \address_gen[22].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[22].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_13 \address_gen[21].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[21].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_12 \address_gen[20].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[20].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_10 \address_gen[19].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[19].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_9 \address_gen[18].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[18].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_8 \address_gen[17].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[17].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_7 \address_gen[16].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[16].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_6 \address_gen[15].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[15].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_5 \address_gen[14].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[14].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_4 \address_gen[13].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[13].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_3 \address_gen[12].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[12].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_2 \address_gen[11].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[11].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_1 \address_gen[10].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[10].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_24 \address_gen[9].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[9].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_23 \address_gen[8].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[8].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_22 \address_gen[7].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[7].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_21 \address_gen[6].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[6].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_20 \address_gen[5].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[5].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_19 \address_gen[4].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[4].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_18 \address_gen[3].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[3].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_17 \address_gen[2].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[2].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc_11 \address_gen[1].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[1].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

system_hps_sdram_p0_acv_ldc \address_gen[0].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[0].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_clk_phase_select \clock_gen[0].clk_phase_select_dqs (
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\clock_gen[0].leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(\mem_ck_source[0] ));
defparam \clock_gen[0].clk_phase_select_dqs .invert_phase = "false";
defparam \clock_gen[0].clk_phase_select_dqs .phase_setting = 0;
defparam \clock_gen[0].clk_phase_select_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].clk_phase_select_dqs .use_dqs_input = "false";
defparam \clock_gen[0].clk_phase_select_dqs .use_phasectrlin = "false";

cyclonev_leveling_delay_chain \clock_gen[0].leveling_delay_chain_dqs (
	.clkin(afi_clk),
	.delayctrlin({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.clkout(\clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ));
defparam \clock_gen[0].leveling_delay_chain_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_delay_increment = 10;
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_intrinsic_delay = 175;

endmodule

module system_altddio_out_1 (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
inout 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_ddio_out_uqe auto_generated(
	.dataout({dataout[0]}),
	.datain_h({datain_h[0]}),
	.datain_l({datain_l[0]}),
	.outclock(outclock));

endmodule

module system_ddio_out_uqe (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
output 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "none";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_acv_ldc (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_1 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_2 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_3 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_4 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_5 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_6 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_7 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_8 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_9 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_10 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_11 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_12 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_13 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_14 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_15 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_16 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_17 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_18 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_19 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_20 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_21 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_22 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_23 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_acv_ldc_24 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_p0_clock_pair_generator (
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	datain)/* synthesis synthesis_greybox=0 */;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	[0:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(datain[0]),
	.oein(gnd),
	.dtcin(gnd),
	.o(wire_pseudo_diffa_o_0),
	.obar(wire_pseudo_diffa_obar_0),
	.oeout(wire_pseudo_diffa_oeout_0),
	.oebout(wire_pseudo_diffa_oebout_0),
	.dtc(),
	.dtcbar());

endmodule

module system_hps_sdram_p0_generic_ddio (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[6].fr_data_lo ;
wire \acblock[6].fr_data_hi ;
wire \acblock[7].fr_data_lo ;
wire \acblock[7].fr_data_hi ;
wire \acblock[8].fr_data_lo ;
wire \acblock[8].fr_data_hi ;
wire \acblock[9].fr_data_lo ;
wire \acblock[9].fr_data_hi ;
wire \acblock[10].fr_data_lo ;
wire \acblock[10].fr_data_hi ;
wire \acblock[11].fr_data_lo ;
wire \acblock[11].fr_data_hi ;
wire \acblock[12].fr_data_lo ;
wire \acblock[12].fr_data_hi ;
wire \acblock[13].fr_data_lo ;
wire \acblock[13].fr_data_hi ;
wire \acblock[14].fr_data_lo ;
wire \acblock[14].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].ddio_out (
	.datainlo(\acblock[6].fr_data_lo ),
	.datainhi(\acblock[6].fr_data_hi ),
	.clkhi(clk_fr[6]),
	.clklo(clk_fr[6]),
	.muxsel(clk_fr[6]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[6]),
	.dfflo(),
	.dffhi());
defparam \acblock[6].ddio_out .async_mode = "none";
defparam \acblock[6].ddio_out .half_rate_mode = "false";
defparam \acblock[6].ddio_out .power_up = "low";
defparam \acblock[6].ddio_out .sync_mode = "none";
defparam \acblock[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].ddio_out (
	.datainlo(\acblock[7].fr_data_lo ),
	.datainhi(\acblock[7].fr_data_hi ),
	.clkhi(clk_fr[7]),
	.clklo(clk_fr[7]),
	.muxsel(clk_fr[7]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[7]),
	.dfflo(),
	.dffhi());
defparam \acblock[7].ddio_out .async_mode = "none";
defparam \acblock[7].ddio_out .half_rate_mode = "false";
defparam \acblock[7].ddio_out .power_up = "low";
defparam \acblock[7].ddio_out .sync_mode = "none";
defparam \acblock[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].ddio_out (
	.datainlo(\acblock[8].fr_data_lo ),
	.datainhi(\acblock[8].fr_data_hi ),
	.clkhi(clk_fr[8]),
	.clklo(clk_fr[8]),
	.muxsel(clk_fr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[8]),
	.dfflo(),
	.dffhi());
defparam \acblock[8].ddio_out .async_mode = "none";
defparam \acblock[8].ddio_out .half_rate_mode = "false";
defparam \acblock[8].ddio_out .power_up = "low";
defparam \acblock[8].ddio_out .sync_mode = "none";
defparam \acblock[8].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].ddio_out (
	.datainlo(\acblock[9].fr_data_lo ),
	.datainhi(\acblock[9].fr_data_hi ),
	.clkhi(clk_fr[9]),
	.clklo(clk_fr[9]),
	.muxsel(clk_fr[9]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[9]),
	.dfflo(),
	.dffhi());
defparam \acblock[9].ddio_out .async_mode = "none";
defparam \acblock[9].ddio_out .half_rate_mode = "false";
defparam \acblock[9].ddio_out .power_up = "low";
defparam \acblock[9].ddio_out .sync_mode = "none";
defparam \acblock[9].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].ddio_out (
	.datainlo(\acblock[10].fr_data_lo ),
	.datainhi(\acblock[10].fr_data_hi ),
	.clkhi(clk_fr[10]),
	.clklo(clk_fr[10]),
	.muxsel(clk_fr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[10]),
	.dfflo(),
	.dffhi());
defparam \acblock[10].ddio_out .async_mode = "none";
defparam \acblock[10].ddio_out .half_rate_mode = "false";
defparam \acblock[10].ddio_out .power_up = "low";
defparam \acblock[10].ddio_out .sync_mode = "none";
defparam \acblock[10].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].ddio_out (
	.datainlo(\acblock[11].fr_data_lo ),
	.datainhi(\acblock[11].fr_data_hi ),
	.clkhi(clk_fr[11]),
	.clklo(clk_fr[11]),
	.muxsel(clk_fr[11]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[11]),
	.dfflo(),
	.dffhi());
defparam \acblock[11].ddio_out .async_mode = "none";
defparam \acblock[11].ddio_out .half_rate_mode = "false";
defparam \acblock[11].ddio_out .power_up = "low";
defparam \acblock[11].ddio_out .sync_mode = "none";
defparam \acblock[11].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].ddio_out (
	.datainlo(\acblock[12].fr_data_lo ),
	.datainhi(\acblock[12].fr_data_hi ),
	.clkhi(clk_fr[12]),
	.clklo(clk_fr[12]),
	.muxsel(clk_fr[12]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[12]),
	.dfflo(),
	.dffhi());
defparam \acblock[12].ddio_out .async_mode = "none";
defparam \acblock[12].ddio_out .half_rate_mode = "false";
defparam \acblock[12].ddio_out .power_up = "low";
defparam \acblock[12].ddio_out .sync_mode = "none";
defparam \acblock[12].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].ddio_out (
	.datainlo(\acblock[13].fr_data_lo ),
	.datainhi(\acblock[13].fr_data_hi ),
	.clkhi(clk_fr[13]),
	.clklo(clk_fr[13]),
	.muxsel(clk_fr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[13]),
	.dfflo(),
	.dffhi());
defparam \acblock[13].ddio_out .async_mode = "none";
defparam \acblock[13].ddio_out .half_rate_mode = "false";
defparam \acblock[13].ddio_out .power_up = "low";
defparam \acblock[13].ddio_out .sync_mode = "none";
defparam \acblock[13].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].ddio_out (
	.datainlo(\acblock[14].fr_data_lo ),
	.datainhi(\acblock[14].fr_data_hi ),
	.clkhi(clk_fr[14]),
	.clklo(clk_fr[14]),
	.muxsel(clk_fr[14]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[14]),
	.dfflo(),
	.dffhi());
defparam \acblock[14].ddio_out .async_mode = "none";
defparam \acblock[14].ddio_out .half_rate_mode = "false";
defparam \acblock[14].ddio_out .power_up = "low";
defparam \acblock[14].ddio_out .sync_mode = "none";
defparam \acblock[14].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_lo (
	.datainlo(datain[27]),
	.datainhi(datain[25]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_lo .async_mode = "none";
defparam \acblock[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_lo .power_up = "low";
defparam \acblock[6].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_hi (
	.datainlo(datain[26]),
	.datainhi(datain[24]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_hi .async_mode = "none";
defparam \acblock[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_hi .power_up = "low";
defparam \acblock[6].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_lo (
	.datainlo(datain[31]),
	.datainhi(datain[29]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_lo .async_mode = "none";
defparam \acblock[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_lo .power_up = "low";
defparam \acblock[7].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_hi (
	.datainlo(datain[30]),
	.datainhi(datain[28]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_hi .async_mode = "none";
defparam \acblock[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_hi .power_up = "low";
defparam \acblock[7].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_lo (
	.datainlo(datain[35]),
	.datainhi(datain[33]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_lo .async_mode = "none";
defparam \acblock[8].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_lo .power_up = "low";
defparam \acblock[8].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[8].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_hi (
	.datainlo(datain[34]),
	.datainhi(datain[32]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_hi .async_mode = "none";
defparam \acblock[8].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_hi .power_up = "low";
defparam \acblock[8].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[8].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_lo (
	.datainlo(datain[39]),
	.datainhi(datain[37]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_lo .async_mode = "none";
defparam \acblock[9].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_lo .power_up = "low";
defparam \acblock[9].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[9].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_hi (
	.datainlo(datain[38]),
	.datainhi(datain[36]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_hi .async_mode = "none";
defparam \acblock[9].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_hi .power_up = "low";
defparam \acblock[9].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[9].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_lo (
	.datainlo(datain[43]),
	.datainhi(datain[41]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_lo .async_mode = "none";
defparam \acblock[10].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_lo .power_up = "low";
defparam \acblock[10].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[10].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_hi (
	.datainlo(datain[42]),
	.datainhi(datain[40]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_hi .async_mode = "none";
defparam \acblock[10].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_hi .power_up = "low";
defparam \acblock[10].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[10].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_lo (
	.datainlo(datain[47]),
	.datainhi(datain[45]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_lo .async_mode = "none";
defparam \acblock[11].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_lo .power_up = "low";
defparam \acblock[11].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[11].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_hi (
	.datainlo(datain[46]),
	.datainhi(datain[44]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_hi .async_mode = "none";
defparam \acblock[11].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_hi .power_up = "low";
defparam \acblock[11].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[11].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_lo (
	.datainlo(datain[51]),
	.datainhi(datain[49]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_lo .async_mode = "none";
defparam \acblock[12].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_lo .power_up = "low";
defparam \acblock[12].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[12].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_hi (
	.datainlo(datain[50]),
	.datainhi(datain[48]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_hi .async_mode = "none";
defparam \acblock[12].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_hi .power_up = "low";
defparam \acblock[12].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[12].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_lo (
	.datainlo(datain[55]),
	.datainhi(datain[53]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_lo .async_mode = "none";
defparam \acblock[13].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_lo .power_up = "low";
defparam \acblock[13].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[13].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_hi (
	.datainlo(datain[54]),
	.datainhi(datain[52]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_hi .async_mode = "none";
defparam \acblock[13].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_hi .power_up = "low";
defparam \acblock[13].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[13].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_lo (
	.datainlo(datain[59]),
	.datainhi(datain[57]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_lo .async_mode = "none";
defparam \acblock[14].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_lo .power_up = "low";
defparam \acblock[14].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[14].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_hi (
	.datainlo(datain[58]),
	.datainhi(datain[56]),
	.clkhi(clk_hr[10]),
	.clklo(clk_hr[10]),
	.muxsel(clk_hr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_hi .async_mode = "none";
defparam \acblock[14].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_hi .power_up = "low";
defparam \acblock[14].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[14].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_generic_ddio_1 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_generic_ddio_2 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_generic_ddio_3 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_altdqdqs (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.write_strobe_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_3,phy_ddio_dmdout_2,phy_ddio_dmdout_1,phy_ddio_dmdout_0}),
	.write_data_in({phy_ddio_dqdout_31,phy_ddio_dqdout_30,phy_ddio_dqdout_29,phy_ddio_dqdout_28,phy_ddio_dqdout_27,phy_ddio_dqdout_26,phy_ddio_dqdout_25,phy_ddio_dqdout_24,phy_ddio_dqdout_23,phy_ddio_dqdout_22,phy_ddio_dqdout_21,phy_ddio_dqdout_20,phy_ddio_dqdout_19,phy_ddio_dqdout_18,
phy_ddio_dqdout_17,phy_ddio_dqdout_16,phy_ddio_dqdout_15,phy_ddio_dqdout_14,phy_ddio_dqdout_13,phy_ddio_dqdout_12,phy_ddio_dqdout_11,phy_ddio_dqdout_10,phy_ddio_dqdout_9,phy_ddio_dqdout_8,phy_ddio_dqdout_7,phy_ddio_dqdout_6,phy_ddio_dqdout_5,phy_ddio_dqdout_4,
phy_ddio_dqdout_3,phy_ddio_dqdout_2,phy_ddio_dqdout_1,phy_ddio_dqdout_0}),
	.write_oe_in({phy_ddio_dqoe_15,phy_ddio_dqoe_14,phy_ddio_dqoe_13,phy_ddio_dqoe_12,phy_ddio_dqoe_11,phy_ddio_dqoe_10,phy_ddio_dqoe_9,phy_ddio_dqoe_8,phy_ddio_dqoe_7,phy_ddio_dqoe_6,phy_ddio_dqoe_5,phy_ddio_dqoe_4,phy_ddio_dqoe_3,phy_ddio_dqoe_2,phy_ddio_dqoe_1,phy_ddio_dqoe_0}),
	.write_strobe({phy_ddio_dqs_dout_3,phy_ddio_dqs_dout_2,phy_ddio_dqs_dout_1,phy_ddio_dqs_dout_0}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_0),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_0),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_1,phy_ddio_dqslogic_incrdataen_0}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_1,phy_ddio_dqslogic_incwrptr_0}),
	.oct_ena_in({phy_ddio_dqslogic_oct_1,phy_ddio_dqslogic_oct_0}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_4,phy_ddio_dqslogic_readlatency_3,phy_ddio_dqslogic_readlatency_2,phy_ddio_dqslogic_readlatency_1,phy_ddio_dqslogic_readlatency_0}),
	.output_strobe_ena({phy_ddio_dqs_oe_1,phy_ddio_dqs_oe_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	write_strobe_clock_in,
	hr_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	write_strobe_clock_in;
input 	hr_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(write_strobe_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(write_strobe_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_altdqdqs_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.write_strobe_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_7,phy_ddio_dmdout_6,phy_ddio_dmdout_5,phy_ddio_dmdout_4}),
	.write_data_in({phy_ddio_dqdout_67,phy_ddio_dqdout_66,phy_ddio_dqdout_65,phy_ddio_dqdout_64,phy_ddio_dqdout_63,phy_ddio_dqdout_62,phy_ddio_dqdout_61,phy_ddio_dqdout_60,phy_ddio_dqdout_59,phy_ddio_dqdout_58,phy_ddio_dqdout_57,phy_ddio_dqdout_56,phy_ddio_dqdout_55,phy_ddio_dqdout_54,
phy_ddio_dqdout_53,phy_ddio_dqdout_52,phy_ddio_dqdout_51,phy_ddio_dqdout_50,phy_ddio_dqdout_49,phy_ddio_dqdout_48,phy_ddio_dqdout_47,phy_ddio_dqdout_46,phy_ddio_dqdout_45,phy_ddio_dqdout_44,phy_ddio_dqdout_43,phy_ddio_dqdout_42,phy_ddio_dqdout_41,phy_ddio_dqdout_40,
phy_ddio_dqdout_39,phy_ddio_dqdout_38,phy_ddio_dqdout_37,phy_ddio_dqdout_36}),
	.write_oe_in({phy_ddio_dqoe_33,phy_ddio_dqoe_32,phy_ddio_dqoe_31,phy_ddio_dqoe_30,phy_ddio_dqoe_29,phy_ddio_dqoe_28,phy_ddio_dqoe_27,phy_ddio_dqoe_26,phy_ddio_dqoe_25,phy_ddio_dqoe_24,phy_ddio_dqoe_23,phy_ddio_dqoe_22,phy_ddio_dqoe_21,phy_ddio_dqoe_20,phy_ddio_dqoe_19,phy_ddio_dqoe_18}),
	.write_strobe({phy_ddio_dqs_dout_7,phy_ddio_dqs_dout_6,phy_ddio_dqs_dout_5,phy_ddio_dqs_dout_4}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_1),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_1),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_3,phy_ddio_dqslogic_incrdataen_2}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_3,phy_ddio_dqslogic_incwrptr_2}),
	.oct_ena_in({phy_ddio_dqslogic_oct_3,phy_ddio_dqslogic_oct_2}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_9,phy_ddio_dqslogic_readlatency_8,phy_ddio_dqslogic_readlatency_7,phy_ddio_dqslogic_readlatency_6,phy_ddio_dqslogic_readlatency_5}),
	.output_strobe_ena({phy_ddio_dqs_oe_3,phy_ddio_dqs_oe_2}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	write_strobe_clock_in,
	hr_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	write_strobe_clock_in;
input 	hr_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(write_strobe_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(write_strobe_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_altdqdqs_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.write_strobe_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_11,phy_ddio_dmdout_10,phy_ddio_dmdout_9,phy_ddio_dmdout_8}),
	.write_data_in({phy_ddio_dqdout_103,phy_ddio_dqdout_102,phy_ddio_dqdout_101,phy_ddio_dqdout_100,phy_ddio_dqdout_99,phy_ddio_dqdout_98,phy_ddio_dqdout_97,phy_ddio_dqdout_96,phy_ddio_dqdout_95,phy_ddio_dqdout_94,phy_ddio_dqdout_93,phy_ddio_dqdout_92,phy_ddio_dqdout_91,phy_ddio_dqdout_90,
phy_ddio_dqdout_89,phy_ddio_dqdout_88,phy_ddio_dqdout_87,phy_ddio_dqdout_86,phy_ddio_dqdout_85,phy_ddio_dqdout_84,phy_ddio_dqdout_83,phy_ddio_dqdout_82,phy_ddio_dqdout_81,phy_ddio_dqdout_80,phy_ddio_dqdout_79,phy_ddio_dqdout_78,phy_ddio_dqdout_77,phy_ddio_dqdout_76,
phy_ddio_dqdout_75,phy_ddio_dqdout_74,phy_ddio_dqdout_73,phy_ddio_dqdout_72}),
	.write_oe_in({phy_ddio_dqoe_51,phy_ddio_dqoe_50,phy_ddio_dqoe_49,phy_ddio_dqoe_48,phy_ddio_dqoe_47,phy_ddio_dqoe_46,phy_ddio_dqoe_45,phy_ddio_dqoe_44,phy_ddio_dqoe_43,phy_ddio_dqoe_42,phy_ddio_dqoe_41,phy_ddio_dqoe_40,phy_ddio_dqoe_39,phy_ddio_dqoe_38,phy_ddio_dqoe_37,phy_ddio_dqoe_36}),
	.write_strobe({phy_ddio_dqs_dout_11,phy_ddio_dqs_dout_10,phy_ddio_dqs_dout_9,phy_ddio_dqs_dout_8}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_2),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_2),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_5,phy_ddio_dqslogic_incrdataen_4}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_5,phy_ddio_dqslogic_incwrptr_4}),
	.oct_ena_in({phy_ddio_dqslogic_oct_5,phy_ddio_dqslogic_oct_4}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_14,phy_ddio_dqslogic_readlatency_13,phy_ddio_dqslogic_readlatency_12,phy_ddio_dqslogic_readlatency_11,phy_ddio_dqslogic_readlatency_10}),
	.output_strobe_ena({phy_ddio_dqs_oe_5,phy_ddio_dqs_oe_4}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	write_strobe_clock_in,
	hr_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	write_strobe_clock_in;
input 	hr_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(write_strobe_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(write_strobe_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_altdqdqs_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.write_strobe_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_15,phy_ddio_dmdout_14,phy_ddio_dmdout_13,phy_ddio_dmdout_12}),
	.write_data_in({phy_ddio_dqdout_139,phy_ddio_dqdout_138,phy_ddio_dqdout_137,phy_ddio_dqdout_136,phy_ddio_dqdout_135,phy_ddio_dqdout_134,phy_ddio_dqdout_133,phy_ddio_dqdout_132,phy_ddio_dqdout_131,phy_ddio_dqdout_130,phy_ddio_dqdout_129,phy_ddio_dqdout_128,phy_ddio_dqdout_127,
phy_ddio_dqdout_126,phy_ddio_dqdout_125,phy_ddio_dqdout_124,phy_ddio_dqdout_123,phy_ddio_dqdout_122,phy_ddio_dqdout_121,phy_ddio_dqdout_120,phy_ddio_dqdout_119,phy_ddio_dqdout_118,phy_ddio_dqdout_117,phy_ddio_dqdout_116,phy_ddio_dqdout_115,phy_ddio_dqdout_114,
phy_ddio_dqdout_113,phy_ddio_dqdout_112,phy_ddio_dqdout_111,phy_ddio_dqdout_110,phy_ddio_dqdout_109,phy_ddio_dqdout_108}),
	.write_oe_in({phy_ddio_dqoe_69,phy_ddio_dqoe_68,phy_ddio_dqoe_67,phy_ddio_dqoe_66,phy_ddio_dqoe_65,phy_ddio_dqoe_64,phy_ddio_dqoe_63,phy_ddio_dqoe_62,phy_ddio_dqoe_61,phy_ddio_dqoe_60,phy_ddio_dqoe_59,phy_ddio_dqoe_58,phy_ddio_dqoe_57,phy_ddio_dqoe_56,phy_ddio_dqoe_55,phy_ddio_dqoe_54}),
	.write_strobe({phy_ddio_dqs_dout_15,phy_ddio_dqs_dout_14,phy_ddio_dqs_dout_13,phy_ddio_dqs_dout_12}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_3),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_3),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_7,phy_ddio_dqslogic_incrdataen_6}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_7,phy_ddio_dqslogic_incwrptr_6}),
	.oct_ena_in({phy_ddio_dqslogic_oct_7,phy_ddio_dqslogic_oct_6}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_19,phy_ddio_dqslogic_readlatency_18,phy_ddio_dqslogic_readlatency_17,phy_ddio_dqslogic_readlatency_16,phy_ddio_dqslogic_readlatency_15}),
	.output_strobe_ena({phy_ddio_dqs_oe_7,phy_ddio_dqs_oe_6}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	write_strobe_clock_in,
	hr_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	write_strobe_clock_in;
input 	hr_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(write_strobe_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(write_strobe_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(write_strobe_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module system_hps_sdram_p0_acv_ldc_25 (
	pll_hr_clk,
	pll_dqs_clk,
	adc_clk,
	avl_clk,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_hr_clk;
input 	pll_dqs_clk;
output 	adc_clk;
output 	avl_clk;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;

assign adc_clk = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

assign avl_clk = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_hr_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(pll_hr_clk),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

endmodule

module system_hps_sdram_pll (
	afi_half_clk,
	pll_write_clk_pre_phy_clk)/* synthesis synthesis_greybox=0 */;
output 	afi_half_clk;
output 	pll_write_clk_pre_phy_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_out[2] ;
wire \clk_out[3] ;

wire [3:0] pll_CLK_OUT_bus;

assign afi_half_clk = pll_CLK_OUT_bus[0];
assign pll_write_clk_pre_phy_clk = pll_CLK_OUT_bus[1];
assign \clk_out[2]  = pll_CLK_OUT_bus[2];
assign \clk_out[3]  = pll_CLK_OUT_bus[3];

cyclonev_hps_sdram_pll pll(
	.ref_clk(gnd),
	.clk_out(pll_CLK_OUT_bus));

endmodule

module system_system_mm_interconnect_0 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	in_data_reg_0,
	int_nxt_addr_reg_dly_1,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	sink1_ready,
	hps_0_h2f_lw_axi_master_awready,
	src0_valid,
	source_endofpacket,
	src1_valid,
	hps_0_h2f_lw_axi_master_wready,
	mem_70_0,
	mem_71_0,
	mem_72_0,
	mem_73_0,
	mem_74_0,
	mem_75_0,
	mem_76_0,
	mem_77_0,
	mem_78_0,
	mem_79_0,
	mem_80_0,
	mem_81_0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	ShiftLeft2,
	ShiftLeft21,
	ShiftLeft22,
	ShiftLeft23,
	ShiftLeft24,
	ShiftLeft25,
	ShiftLeft26,
	ShiftLeft27,
	ShiftLeft28,
	ShiftLeft29,
	ShiftLeft210,
	ShiftLeft211,
	ShiftLeft212,
	ShiftLeft213,
	ShiftLeft214,
	ShiftLeft215,
	m0_write,
	source0_data_16,
	source0_data_17,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_1;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	sink1_ready;
output 	hps_0_h2f_lw_axi_master_awready;
output 	src0_valid;
output 	source_endofpacket;
output 	src1_valid;
output 	hps_0_h2f_lw_axi_master_wready;
output 	mem_70_0;
output 	mem_71_0;
output 	mem_72_0;
output 	mem_73_0;
output 	mem_74_0;
output 	mem_75_0;
output 	mem_76_0;
output 	mem_77_0;
output 	mem_78_0;
output 	mem_79_0;
output 	mem_80_0;
output 	mem_81_0;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	ShiftLeft2;
output 	ShiftLeft21;
output 	ShiftLeft22;
output 	ShiftLeft23;
output 	ShiftLeft24;
output 	ShiftLeft25;
output 	ShiftLeft26;
output 	ShiftLeft27;
output 	ShiftLeft28;
output 	ShiftLeft29;
output 	ShiftLeft210;
output 	ShiftLeft211;
output 	ShiftLeft212;
output 	ShiftLeft213;
output 	ShiftLeft214;
output 	ShiftLeft215;
output 	m0_write;
output 	source0_data_16;
output 	source0_data_17;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_0_h2f_lw_axi_master_agent|Add4~1_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~1_sumout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[1]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[0]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~5_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~5_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~9_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~9_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~13_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~13_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~17_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~17_sumout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ;
wire \ram_s1_cmd_width_adapter|out_data[49]~36_combout ;
wire \cmd_mux|src_data[66]~24_combout ;
wire \ram_s1_rsp_width_adapter|always10~1_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \cmd_mux|saved_grant[0]~q ;
wire \cmd_mux|src_data[78]~combout ;
wire \cmd_mux|src_data[79]~combout ;
wire \cmd_mux|src_data[77]~combout ;
wire \ram_s1_cmd_width_adapter|in_ready~0_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \ram_s1_agent|WideOr0~combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ;
wire \ram_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ;
wire \cmd_mux|src_valid~0_combout ;
wire \ram_s1_translator|read_latency_shift_reg[0]~q ;
wire \ram_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \ram_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \ram_s1_rsp_width_adapter|out_valid~0_combout ;
wire \ram_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \ram_s1_agent|comb~0_combout ;
wire \ram_s1_agent_rsp_fifo|mem[0][39]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][51]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][50]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][49]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][48]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][47]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][46]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][45]~q ;
wire \ram_s1_agent|uncompressor|last_packet_beat~4_combout ;
wire \ram_s1_agent|uncompressor|source_addr[1]~0_combout ;
wire \ram_s1_agent|uncompressor|source_addr[1]~1_combout ;
wire \ram_s1_agent_rsp_fifo|mem[0][19]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][91]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][59]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][41]~q ;
wire \rsp_demux|src0_valid~0_combout ;
wire \ram_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][10]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][11]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][12]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][13]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][14]~q ;
wire \ram_s1_agent_rdata_fifo|mem[0][15]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[41]~q ;
wire \ram_s1_agent|m0_write~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ;
wire \ram_s1_cmd_width_adapter|use_reg~q ;
wire \cmd_mux|WideOr1~combout ;
wire \ram_s1_cmd_width_adapter|out_endofpacket~1_combout ;
wire \ram_s1_cmd_width_adapter|out_data[59]~0_combout ;
wire \cmd_mux|src_payload~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add1~0_combout ;
wire \cmd_mux|src_payload~3_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add3~0_combout ;
wire \cmd_mux|src_data[70]~3_combout ;
wire \hps_0_h2f_lw_axi_master_agent|sop_enable~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[0]~q ;
wire \ram_s1_cmd_width_adapter|out_data[18]~2_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[1]~q ;
wire \ram_s1_cmd_width_adapter|int_output_sel[0]~1_combout ;
wire \ram_s1_cmd_width_adapter|out_data[17]~3_combout ;
wire \ram_s1_cmd_width_adapter|out_data[16]~4_combout ;
wire \ram_s1_rsp_width_adapter|p1_ready~0_combout ;
wire \ram_s1_agent|uncompressor|sink_ready~0_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[42]~q ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ;
wire \cmd_mux|src_payload~5_combout ;
wire \cmd_mux|src_data[69]~combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[5]~q ;
wire \hps_0_h2f_lw_axi_master_agent|Add6~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add2~0_combout ;
wire \cmd_mux|src_data[68]~combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[4]~q ;
wire \hps_0_h2f_lw_axi_master_agent|Add6~1_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add2~1_combout ;
wire \cmd_mux|src_data[67]~combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[3]~q ;
wire \hps_0_h2f_lw_axi_master_agent|Add2~2_combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[2]~q ;
wire \cmd_mux|src_data[65]~combout ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ;
wire \cmd_mux|src_payload~6_combout ;
wire \ram_s1_cmd_width_adapter|out_data[50]~8_combout ;
wire \ram_s1_cmd_width_adapter|out_data[48]~9_combout ;
wire \ram_s1_cmd_width_adapter|ShiftLeft0~1_combout ;
wire \ram_s1_cmd_width_adapter|out_data[47]~10_combout ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ;
wire \ram_s1_cmd_width_adapter|out_data[47]~12_combout ;
wire \ram_s1_cmd_width_adapter|out_data[51]~13_combout ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ;
wire \cmd_mux|src_payload~7_combout ;
wire \ram_s1_cmd_width_adapter|out_data[51]~15_combout ;
wire \ram_s1_cmd_width_adapter|byte_cnt_reg[1]~q ;
wire \ram_s1_cmd_width_adapter|out_data[46]~16_combout ;
wire \ram_s1_cmd_width_adapter|out_data[46]~17_combout ;
wire \ram_s1_agent|cp_ready~0_combout ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[1]~q ;
wire \ram_s1_rsp_width_adapter|out_valid~1_combout ;
wire \ram_s1_agent_rsp_fifo|mem[0][53]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[70]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[71]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[72]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[73]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[74]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[75]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[76]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[77]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[78]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[79]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[80]~q ;
wire \ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[81]~q ;
wire \ram_s1_cmd_width_adapter|out_data[0]~18_combout ;
wire \cmd_mux|src_payload~8_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add1~1_combout ;
wire \cmd_mux|src_payload~9_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add3~1_combout ;
wire \cmd_mux|src_data[71]~5_combout ;
wire \cmd_mux|src_payload~10_combout ;
wire \hps_0_h2f_lw_axi_master_agent|LessThan12~0_combout ;
wire \cmd_mux|src_payload~11_combout ;
wire \cmd_mux|src_data[72]~8_combout ;
wire \ram_s1_cmd_width_adapter|address_reg[2]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[2]~q ;
wire \cmd_mux|src_data[38]~combout ;
wire \cmd_mux|src_payload~12_combout ;
wire \cmd_mux|src_data[73]~11_combout ;
wire \ram_s1_cmd_width_adapter|address_reg[3]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[3]~q ;
wire \cmd_mux|src_data[39]~combout ;
wire \cmd_mux|src_payload~13_combout ;
wire \cmd_mux|src_payload~14_combout ;
wire \cmd_mux|src_data[74]~13_combout ;
wire \ram_s1_cmd_width_adapter|address_reg[4]~q ;
wire \cmd_mux|src_payload~15_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~0_combout ;
wire \ram_s1_cmd_width_adapter|out_data[1]~19_combout ;
wire \ram_s1_cmd_width_adapter|out_data[2]~20_combout ;
wire \ram_s1_cmd_width_adapter|out_data[3]~21_combout ;
wire \ram_s1_cmd_width_adapter|out_data[4]~22_combout ;
wire \ram_s1_cmd_width_adapter|out_data[5]~23_combout ;
wire \ram_s1_cmd_width_adapter|out_data[6]~24_combout ;
wire \ram_s1_cmd_width_adapter|out_data[7]~25_combout ;
wire \ram_s1_cmd_width_adapter|out_data[8]~26_combout ;
wire \ram_s1_cmd_width_adapter|out_data[9]~27_combout ;
wire \ram_s1_cmd_width_adapter|out_data[10]~28_combout ;
wire \ram_s1_cmd_width_adapter|out_data[11]~29_combout ;
wire \ram_s1_cmd_width_adapter|out_data[12]~30_combout ;
wire \ram_s1_cmd_width_adapter|out_data[13]~31_combout ;
wire \ram_s1_cmd_width_adapter|out_data[14]~32_combout ;
wire \ram_s1_cmd_width_adapter|out_data[15]~33_combout ;
wire \cmd_mux|src_payload[0]~combout ;
wire \cmd_mux|src_data[70]~15_combout ;
wire \ram_s1_cmd_width_adapter|out_data[48]~34_combout ;
wire \ram_s1_cmd_width_adapter|out_data[51]~35_combout ;
wire \cmd_mux|src_data[88]~combout ;
wire \cmd_mux|src_data[89]~combout ;
wire \cmd_mux|src_data[90]~combout ;
wire \cmd_mux|src_data[91]~combout ;
wire \cmd_mux|src_data[92]~combout ;
wire \cmd_mux|src_data[93]~combout ;
wire \cmd_mux|src_data[94]~combout ;
wire \cmd_mux|src_data[95]~combout ;
wire \cmd_mux|src_data[96]~combout ;
wire \cmd_mux|src_data[97]~combout ;
wire \cmd_mux|src_data[98]~combout ;
wire \cmd_mux|src_data[99]~combout ;
wire \cmd_mux|src_data[71]~17_combout ;
wire \cmd_mux|src_data[72]~19_combout ;
wire \cmd_mux|src_data[73]~21_combout ;
wire \cmd_mux|src_payload~17_combout ;
wire \cmd_mux|src_data[74]~23_combout ;
wire \ram_s1_agent_rsp_fifo|mem[0][18]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][52]~q ;
wire \ram_s1_agent|cp_ready~1_combout ;


system_altera_avalon_sc_fifo ram_s1_agent_rdata_fifo(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_10(q_a_10),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\ram_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_94_0(\ram_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_used_01(\ram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.mem_0_0(\ram_s1_agent_rdata_fifo|mem[0][0]~q ),
	.mem_1_0(\ram_s1_agent_rdata_fifo|mem[0][1]~q ),
	.mem_2_0(\ram_s1_agent_rdata_fifo|mem[0][2]~q ),
	.mem_3_0(\ram_s1_agent_rdata_fifo|mem[0][3]~q ),
	.mem_4_0(\ram_s1_agent_rdata_fifo|mem[0][4]~q ),
	.mem_5_0(\ram_s1_agent_rdata_fifo|mem[0][5]~q ),
	.mem_6_0(\ram_s1_agent_rdata_fifo|mem[0][6]~q ),
	.mem_7_0(\ram_s1_agent_rdata_fifo|mem[0][7]~q ),
	.mem_8_0(\ram_s1_agent_rdata_fifo|mem[0][8]~q ),
	.mem_9_0(\ram_s1_agent_rdata_fifo|mem[0][9]~q ),
	.mem_10_0(\ram_s1_agent_rdata_fifo|mem[0][10]~q ),
	.mem_11_0(\ram_s1_agent_rdata_fifo|mem[0][11]~q ),
	.mem_12_0(\ram_s1_agent_rdata_fifo|mem[0][12]~q ),
	.mem_13_0(\ram_s1_agent_rdata_fifo|mem[0][13]~q ),
	.mem_14_0(\ram_s1_agent_rdata_fifo|mem[0][14]~q ),
	.mem_15_0(\ram_s1_agent_rdata_fifo|mem[0][15]~q ),
	.reset(r_sync_rst),
	.p1_ready(\ram_s1_rsp_width_adapter|p1_ready~0_combout ),
	.out_valid(\ram_s1_rsp_width_adapter|out_valid~1_combout ),
	.clk(clk_clk));

system_altera_avalon_sc_fifo_1 ram_s1_agent_rsp_fifo(
	.int_nxt_addr_reg_dly_1(int_nxt_addr_reg_dly_1),
	.out_uncomp_byte_cnt_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[1]~q ),
	.out_uncomp_byte_cnt_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[0]~q ),
	.out_uncomp_byte_cnt_reg_5(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_4(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_burstwrap_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ),
	.out_addr_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ),
	.out_burstwrap_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ),
	.nxt_out_eop(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.in_data_reg_59(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.WideOr0(\ram_s1_agent|WideOr0~combout ),
	.mem_used_1(\ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.nxt_out_eop1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.out_valid_reg(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_94_0(\ram_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_used_0(\ram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_95_0(\ram_s1_agent_rsp_fifo|mem[0][95]~q ),
	.comb(\ram_s1_agent|comb~0_combout ),
	.mem_39_0(\ram_s1_agent_rsp_fifo|mem[0][39]~q ),
	.mem_51_0(\ram_s1_agent_rsp_fifo|mem[0][51]~q ),
	.mem_50_0(\ram_s1_agent_rsp_fifo|mem[0][50]~q ),
	.mem_49_0(\ram_s1_agent_rsp_fifo|mem[0][49]~q ),
	.mem_48_0(\ram_s1_agent_rsp_fifo|mem[0][48]~q ),
	.mem_47_0(\ram_s1_agent_rsp_fifo|mem[0][47]~q ),
	.mem_46_0(\ram_s1_agent_rsp_fifo|mem[0][46]~q ),
	.mem_45_0(\ram_s1_agent_rsp_fifo|mem[0][45]~q ),
	.last_packet_beat(\ram_s1_agent|uncompressor|last_packet_beat~4_combout ),
	.mem_19_0(\ram_s1_agent_rsp_fifo|mem[0][19]~q ),
	.mem_91_0(\ram_s1_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\ram_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\ram_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_59_0(\ram_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_41_0(\ram_s1_agent_rsp_fifo|mem[0][41]~q ),
	.mem_70_0(mem_70_0),
	.mem_71_0(mem_71_0),
	.mem_72_0(mem_72_0),
	.mem_73_0(mem_73_0),
	.mem_74_0(mem_74_0),
	.mem_75_0(mem_75_0),
	.mem_76_0(mem_76_0),
	.mem_77_0(mem_77_0),
	.mem_78_0(mem_78_0),
	.mem_79_0(mem_79_0),
	.mem_80_0(mem_80_0),
	.mem_81_0(mem_81_0),
	.in_data_reg_41(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[41]~q ),
	.m0_write(\ram_s1_agent|m0_write~0_combout ),
	.reset(r_sync_rst),
	.p1_ready(\ram_s1_rsp_width_adapter|p1_ready~0_combout ),
	.sink_ready(\ram_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_42(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[42]~q ),
	.out_byte_cnt_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[1]~q ),
	.out_valid(\ram_s1_rsp_width_adapter|out_valid~1_combout ),
	.mem_53_0(\ram_s1_agent_rsp_fifo|mem[0][53]~q ),
	.in_data_reg_91(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_70(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[70]~q ),
	.in_data_reg_71(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[71]~q ),
	.in_data_reg_72(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[72]~q ),
	.in_data_reg_73(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[73]~q ),
	.in_data_reg_74(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[74]~q ),
	.in_data_reg_75(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[75]~q ),
	.in_data_reg_76(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[76]~q ),
	.in_data_reg_77(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[77]~q ),
	.in_data_reg_78(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[78]~q ),
	.in_data_reg_79(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[79]~q ),
	.in_data_reg_80(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[80]~q ),
	.in_data_reg_81(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[81]~q ),
	.mem_18_0(\ram_s1_agent_rsp_fifo|mem[0][18]~q ),
	.mem_52_0(\ram_s1_agent_rsp_fifo|mem[0][52]~q ),
	.cp_ready(\ram_s1_agent|cp_ready~1_combout ),
	.clk(clk_clk));

system_altera_merlin_slave_agent ram_s1_agent(
	.always10(\ram_s1_rsp_width_adapter|always10~1_combout ),
	.stateST_COMP_TRANS(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_narrow_reg(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr01(\ram_s1_agent|WideOr0~combout ),
	.in_ready_hold(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.out_valid_reg(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\ram_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_94_0(\ram_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_used_01(\ram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.out_valid(\ram_s1_rsp_width_adapter|out_valid~0_combout ),
	.mem_95_0(\ram_s1_agent_rsp_fifo|mem[0][95]~q ),
	.comb(\ram_s1_agent|comb~0_combout ),
	.mem_39_0(\ram_s1_agent_rsp_fifo|mem[0][39]~q ),
	.mem_51_0(\ram_s1_agent_rsp_fifo|mem[0][51]~q ),
	.mem_50_0(\ram_s1_agent_rsp_fifo|mem[0][50]~q ),
	.mem_49_0(\ram_s1_agent_rsp_fifo|mem[0][49]~q ),
	.mem_48_0(\ram_s1_agent_rsp_fifo|mem[0][48]~q ),
	.mem_47_0(\ram_s1_agent_rsp_fifo|mem[0][47]~q ),
	.mem_46_0(\ram_s1_agent_rsp_fifo|mem[0][46]~q ),
	.mem_45_0(\ram_s1_agent_rsp_fifo|mem[0][45]~q ),
	.last_packet_beat(\ram_s1_agent|uncompressor|last_packet_beat~4_combout ),
	.source_addr_1(\ram_s1_agent|uncompressor|source_addr[1]~0_combout ),
	.source_addr_11(\ram_s1_agent|uncompressor|source_addr[1]~1_combout ),
	.mem_19_0(\ram_s1_agent_rsp_fifo|mem[0][19]~q ),
	.mem_59_0(\ram_s1_agent_rsp_fifo|mem[0][59]~q ),
	.source_endofpacket(source_endofpacket),
	.in_data_reg_41(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[41]~q ),
	.m0_write(\ram_s1_agent|m0_write~0_combout ),
	.m0_write1(m0_write),
	.r_sync_rst(r_sync_rst),
	.p1_ready(\ram_s1_rsp_width_adapter|p1_ready~0_combout ),
	.rf_sink_ready(\ram_s1_agent|uncompressor|sink_ready~0_combout ),
	.cp_ready(\ram_s1_agent|cp_ready~0_combout ),
	.out_valid1(\ram_s1_rsp_width_adapter|out_valid~1_combout ),
	.mem_53_0(\ram_s1_agent_rsp_fifo|mem[0][53]~q ),
	.mem_18_0(\ram_s1_agent_rsp_fifo|mem[0][18]~q ),
	.mem_52_0(\ram_s1_agent_rsp_fifo|mem[0][52]~q ),
	.cp_ready1(\ram_s1_agent|cp_ready~1_combout ),
	.clk_clk(clk_clk));

system_altera_merlin_axi_master_ni hps_0_h2f_lw_axi_master_agent(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_0(h2f_lw_AWLEN_0),
	.h2f_lw_AWLEN_1(h2f_lw_AWLEN_1),
	.h2f_lw_AWLEN_2(h2f_lw_AWLEN_2),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.Add4(\hps_0_h2f_lw_axi_master_agent|Add4~1_sumout ),
	.Add5(\hps_0_h2f_lw_axi_master_agent|Add5~1_sumout ),
	.Add41(\hps_0_h2f_lw_axi_master_agent|Add4~5_sumout ),
	.Add51(\hps_0_h2f_lw_axi_master_agent|Add5~5_sumout ),
	.Add42(\hps_0_h2f_lw_axi_master_agent|Add4~9_sumout ),
	.Add52(\hps_0_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add43(\hps_0_h2f_lw_axi_master_agent|Add4~13_sumout ),
	.Add53(\hps_0_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Add44(\hps_0_h2f_lw_axi_master_agent|Add4~17_sumout ),
	.Add54(\hps_0_h2f_lw_axi_master_agent|Add5~17_sumout ),
	.in_ready(\ram_s1_cmd_width_adapter|in_ready~0_combout ),
	.nxt_out_eop(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.nxt_out_eop1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.nxt_in_ready(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready2(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.awready(hps_0_h2f_lw_axi_master_awready),
	.wready(hps_0_h2f_lw_axi_master_wready),
	.write_addr_data_both_valid1(\hps_0_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ),
	.Add1(\hps_0_h2f_lw_axi_master_agent|Add1~0_combout ),
	.src_payload(\cmd_mux|src_payload~3_combout ),
	.Add3(\hps_0_h2f_lw_axi_master_agent|Add3~0_combout ),
	.sop_enable1(\hps_0_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_0(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[0]~q ),
	.address_burst_1(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[1]~q ),
	.write_cp_data_69(\hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.burst_bytecount_5(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.Add6(\hps_0_h2f_lw_axi_master_agent|Add6~0_combout ),
	.Add2(\hps_0_h2f_lw_axi_master_agent|Add2~0_combout ),
	.burst_bytecount_4(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.Add61(\hps_0_h2f_lw_axi_master_agent|Add6~1_combout ),
	.Add21(\hps_0_h2f_lw_axi_master_agent|Add2~1_combout ),
	.burst_bytecount_3(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.Add22(\hps_0_h2f_lw_axi_master_agent|Add2~2_combout ),
	.burst_bytecount_2(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_66(\hps_0_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ),
	.write_cp_data_67(\hps_0_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.write_cp_data_68(\hps_0_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ),
	.Add11(\hps_0_h2f_lw_axi_master_agent|Add1~1_combout ),
	.src_payload1(\cmd_mux|src_payload~9_combout ),
	.Add31(\hps_0_h2f_lw_axi_master_agent|Add3~1_combout ),
	.LessThan12(\hps_0_h2f_lw_axi_master_agent|LessThan12~0_combout ),
	.src_payload2(\cmd_mux|src_payload~11_combout ),
	.address_burst_2(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[2]~q ),
	.address_burst_3(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[3]~q ),
	.src_payload3(\cmd_mux|src_payload~14_combout ),
	.out_data_4(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_payload4(\cmd_mux|src_payload~17_combout ),
	.clk_clk(clk_clk));

system_altera_merlin_slave_translator ram_s1_translator(
	.WideOr0(\ram_s1_agent|WideOr0~combout ),
	.in_ready_hold(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write(\ram_s1_agent|m0_write~0_combout ),
	.reset(r_sync_rst),
	.in_data_reg_42(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[42]~q ),
	.clk(clk_clk));

system_altera_merlin_width_adapter ram_s1_cmd_width_adapter(
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.out_data_49(\ram_s1_cmd_width_adapter|out_data[49]~36_combout ),
	.src_data_66(\cmd_mux|src_data[66]~24_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.in_ready(\ram_s1_cmd_width_adapter|in_ready~0_combout ),
	.nxt_out_eop(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.nxt_out_eop1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.nxt_in_ready(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready2(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.r_sync_rst(r_sync_rst),
	.use_reg1(\ram_s1_cmd_width_adapter|use_reg~q ),
	.WideOr1(\cmd_mux|WideOr1~combout ),
	.out_endofpacket(\ram_s1_cmd_width_adapter|out_endofpacket~1_combout ),
	.out_data_59(\ram_s1_cmd_width_adapter|out_data[59]~0_combout ),
	.sop_enable(\hps_0_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_0(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[0]~q ),
	.out_data_18(\ram_s1_cmd_width_adapter|out_data[18]~2_combout ),
	.address_burst_1(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[1]~q ),
	.int_output_sel_0(\ram_s1_cmd_width_adapter|int_output_sel[0]~1_combout ),
	.out_data_17(\ram_s1_cmd_width_adapter|out_data[17]~3_combout ),
	.out_data_16(\ram_s1_cmd_width_adapter|out_data[16]~4_combout ),
	.write_cp_data_69(\hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.src_payload(\cmd_mux|src_payload~5_combout ),
	.src_data_69(\cmd_mux|src_data[69]~combout ),
	.src_data_68(\cmd_mux|src_data[68]~combout ),
	.Add2(\hps_0_h2f_lw_axi_master_agent|Add2~1_combout ),
	.src_data_67(\cmd_mux|src_data[67]~combout ),
	.src_data_65(\cmd_mux|src_data[65]~combout ),
	.write_cp_data_66(\hps_0_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ),
	.src_payload1(\cmd_mux|src_payload~6_combout ),
	.out_data_50(\ram_s1_cmd_width_adapter|out_data[50]~8_combout ),
	.out_data_48(\ram_s1_cmd_width_adapter|out_data[48]~9_combout ),
	.ShiftLeft0(\ram_s1_cmd_width_adapter|ShiftLeft0~1_combout ),
	.out_data_47(\ram_s1_cmd_width_adapter|out_data[47]~10_combout ),
	.write_cp_data_67(\hps_0_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.out_data_471(\ram_s1_cmd_width_adapter|out_data[47]~12_combout ),
	.out_data_51(\ram_s1_cmd_width_adapter|out_data[51]~13_combout ),
	.write_cp_data_68(\hps_0_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ),
	.src_payload2(\cmd_mux|src_payload~7_combout ),
	.out_data_511(\ram_s1_cmd_width_adapter|out_data[51]~15_combout ),
	.byte_cnt_reg_1(\ram_s1_cmd_width_adapter|byte_cnt_reg[1]~q ),
	.out_data_46(\ram_s1_cmd_width_adapter|out_data[46]~16_combout ),
	.out_data_461(\ram_s1_cmd_width_adapter|out_data[46]~17_combout ),
	.out_data_0(\ram_s1_cmd_width_adapter|out_data[0]~18_combout ),
	.address_reg_2(\ram_s1_cmd_width_adapter|address_reg[2]~q ),
	.src_data_38(\cmd_mux|src_data[38]~combout ),
	.address_reg_3(\ram_s1_cmd_width_adapter|address_reg[3]~q ),
	.src_data_39(\cmd_mux|src_data[39]~combout ),
	.address_reg_4(\ram_s1_cmd_width_adapter|address_reg[4]~q ),
	.src_payload3(\cmd_mux|src_payload~15_combout ),
	.out_data_4(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~0_combout ),
	.out_data_1(\ram_s1_cmd_width_adapter|out_data[1]~19_combout ),
	.out_data_2(\ram_s1_cmd_width_adapter|out_data[2]~20_combout ),
	.out_data_3(\ram_s1_cmd_width_adapter|out_data[3]~21_combout ),
	.out_data_41(\ram_s1_cmd_width_adapter|out_data[4]~22_combout ),
	.out_data_5(\ram_s1_cmd_width_adapter|out_data[5]~23_combout ),
	.out_data_6(\ram_s1_cmd_width_adapter|out_data[6]~24_combout ),
	.out_data_7(\ram_s1_cmd_width_adapter|out_data[7]~25_combout ),
	.out_data_8(\ram_s1_cmd_width_adapter|out_data[8]~26_combout ),
	.out_data_9(\ram_s1_cmd_width_adapter|out_data[9]~27_combout ),
	.out_data_10(\ram_s1_cmd_width_adapter|out_data[10]~28_combout ),
	.out_data_11(\ram_s1_cmd_width_adapter|out_data[11]~29_combout ),
	.out_data_12(\ram_s1_cmd_width_adapter|out_data[12]~30_combout ),
	.out_data_13(\ram_s1_cmd_width_adapter|out_data[13]~31_combout ),
	.out_data_14(\ram_s1_cmd_width_adapter|out_data[14]~32_combout ),
	.out_data_15(\ram_s1_cmd_width_adapter|out_data[15]~33_combout ),
	.in_endofpacket(\cmd_mux|src_payload[0]~combout ),
	.out_data_481(\ram_s1_cmd_width_adapter|out_data[48]~34_combout ),
	.out_data_512(\ram_s1_cmd_width_adapter|out_data[51]~35_combout ),
	.clk_clk(clk_clk));

system_altera_merlin_width_adapter_1 ram_s1_rsp_width_adapter(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_10(q_a_10),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.always10(\ram_s1_rsp_width_adapter|always10~1_combout ),
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\ram_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_94_0(\ram_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_used_01(\ram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.out_valid(\ram_s1_rsp_width_adapter|out_valid~0_combout ),
	.mem_95_0(\ram_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_39_0(\ram_s1_agent_rsp_fifo|mem[0][39]~q ),
	.last_packet_beat(\ram_s1_agent|uncompressor|last_packet_beat~4_combout ),
	.source_addr_1(\ram_s1_agent|uncompressor|source_addr[1]~0_combout ),
	.source_addr_11(\ram_s1_agent|uncompressor|source_addr[1]~1_combout ),
	.mem_19_0(\ram_s1_agent_rsp_fifo|mem[0][19]~q ),
	.mem_91_0(\ram_s1_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\ram_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\ram_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_59_0(\ram_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_41_0(\ram_s1_agent_rsp_fifo|mem[0][41]~q ),
	.mem_0_0(\ram_s1_agent_rdata_fifo|mem[0][0]~q ),
	.out_data_0(out_data_0),
	.mem_1_0(\ram_s1_agent_rdata_fifo|mem[0][1]~q ),
	.out_data_1(out_data_1),
	.mem_2_0(\ram_s1_agent_rdata_fifo|mem[0][2]~q ),
	.out_data_2(out_data_2),
	.mem_3_0(\ram_s1_agent_rdata_fifo|mem[0][3]~q ),
	.out_data_3(out_data_3),
	.mem_4_0(\ram_s1_agent_rdata_fifo|mem[0][4]~q ),
	.out_data_4(out_data_4),
	.mem_5_0(\ram_s1_agent_rdata_fifo|mem[0][5]~q ),
	.out_data_5(out_data_5),
	.mem_6_0(\ram_s1_agent_rdata_fifo|mem[0][6]~q ),
	.out_data_6(out_data_6),
	.mem_7_0(\ram_s1_agent_rdata_fifo|mem[0][7]~q ),
	.out_data_7(out_data_7),
	.mem_8_0(\ram_s1_agent_rdata_fifo|mem[0][8]~q ),
	.out_data_8(out_data_8),
	.mem_9_0(\ram_s1_agent_rdata_fifo|mem[0][9]~q ),
	.out_data_9(out_data_9),
	.mem_10_0(\ram_s1_agent_rdata_fifo|mem[0][10]~q ),
	.out_data_10(out_data_10),
	.mem_11_0(\ram_s1_agent_rdata_fifo|mem[0][11]~q ),
	.out_data_11(out_data_11),
	.mem_12_0(\ram_s1_agent_rdata_fifo|mem[0][12]~q ),
	.out_data_12(out_data_12),
	.mem_13_0(\ram_s1_agent_rdata_fifo|mem[0][13]~q ),
	.out_data_13(out_data_13),
	.mem_14_0(\ram_s1_agent_rdata_fifo|mem[0][14]~q ),
	.out_data_14(out_data_14),
	.mem_15_0(\ram_s1_agent_rdata_fifo|mem[0][15]~q ),
	.out_data_15(out_data_15),
	.ShiftLeft2(ShiftLeft2),
	.ShiftLeft21(ShiftLeft21),
	.ShiftLeft22(ShiftLeft22),
	.ShiftLeft23(ShiftLeft23),
	.ShiftLeft24(ShiftLeft24),
	.ShiftLeft25(ShiftLeft25),
	.ShiftLeft26(ShiftLeft26),
	.ShiftLeft27(ShiftLeft27),
	.ShiftLeft28(ShiftLeft28),
	.ShiftLeft29(ShiftLeft29),
	.ShiftLeft210(ShiftLeft210),
	.ShiftLeft211(ShiftLeft211),
	.ShiftLeft212(ShiftLeft212),
	.ShiftLeft213(ShiftLeft213),
	.ShiftLeft214(ShiftLeft214),
	.ShiftLeft215(ShiftLeft215),
	.r_sync_rst(r_sync_rst),
	.p1_ready(\ram_s1_rsp_width_adapter|p1_ready~0_combout ),
	.out_valid1(\ram_s1_rsp_width_adapter|out_valid~1_combout ),
	.clk_clk(clk_clk));

system_system_mm_interconnect_0_rsp_demux rsp_demux(
	.always10(\ram_s1_rsp_width_adapter|always10~1_combout ),
	.out_valid(\ram_s1_rsp_width_adapter|out_valid~0_combout ),
	.mem_95_0(\ram_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_39_0(\ram_s1_agent_rsp_fifo|mem[0][39]~q ),
	.last_packet_beat(\ram_s1_agent|uncompressor|last_packet_beat~4_combout ),
	.mem_41_0(\ram_s1_agent_rsp_fifo|mem[0][41]~q ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.src0_valid1(src0_valid),
	.src1_valid(src1_valid));

system_system_mm_interconnect_0_cmd_mux cmd_mux(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWLEN_0(h2f_lw_AWLEN_0),
	.h2f_lw_AWLEN_1(h2f_lw_AWLEN_1),
	.h2f_lw_AWLEN_2(h2f_lw_AWLEN_2),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.Add4(\hps_0_h2f_lw_axi_master_agent|Add4~1_sumout ),
	.Add5(\hps_0_h2f_lw_axi_master_agent|Add5~1_sumout ),
	.Add41(\hps_0_h2f_lw_axi_master_agent|Add4~5_sumout ),
	.Add51(\hps_0_h2f_lw_axi_master_agent|Add5~5_sumout ),
	.Add42(\hps_0_h2f_lw_axi_master_agent|Add4~9_sumout ),
	.Add52(\hps_0_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add43(\hps_0_h2f_lw_axi_master_agent|Add4~13_sumout ),
	.Add53(\hps_0_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Add44(\hps_0_h2f_lw_axi_master_agent|Add4~17_sumout ),
	.Add54(\hps_0_h2f_lw_axi_master_agent|Add5~17_sumout ),
	.src_data_66(\cmd_mux|src_data[66]~24_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.in_ready(\ram_s1_cmd_width_adapter|in_ready~0_combout ),
	.nxt_out_eop(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.nxt_out_eop1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.nxt_in_ready(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.sink1_ready1(sink1_ready),
	.nxt_in_ready2(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.write_addr_data_both_valid(\hps_0_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ),
	.r_sync_rst(r_sync_rst),
	.WideOr11(\cmd_mux|WideOr1~combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.Add1(\hps_0_h2f_lw_axi_master_agent|Add1~0_combout ),
	.src_payload1(\cmd_mux|src_payload~3_combout ),
	.Add3(\hps_0_h2f_lw_axi_master_agent|Add3~0_combout ),
	.src_data_70(\cmd_mux|src_data[70]~3_combout ),
	.sop_enable(\hps_0_h2f_lw_axi_master_agent|sop_enable~q ),
	.write_cp_data_69(\hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.src_payload2(\cmd_mux|src_payload~5_combout ),
	.src_data_69(\cmd_mux|src_data[69]~combout ),
	.burst_bytecount_5(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.Add6(\hps_0_h2f_lw_axi_master_agent|Add6~0_combout ),
	.Add2(\hps_0_h2f_lw_axi_master_agent|Add2~0_combout ),
	.src_data_68(\cmd_mux|src_data[68]~combout ),
	.burst_bytecount_4(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.Add61(\hps_0_h2f_lw_axi_master_agent|Add6~1_combout ),
	.Add21(\hps_0_h2f_lw_axi_master_agent|Add2~1_combout ),
	.src_data_67(\cmd_mux|src_data[67]~combout ),
	.burst_bytecount_3(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.Add22(\hps_0_h2f_lw_axi_master_agent|Add2~2_combout ),
	.burst_bytecount_2(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.src_data_65(\cmd_mux|src_data[65]~combout ),
	.src_payload3(\cmd_mux|src_payload~6_combout ),
	.src_payload4(\cmd_mux|src_payload~7_combout ),
	.src_payload5(\cmd_mux|src_payload~8_combout ),
	.Add11(\hps_0_h2f_lw_axi_master_agent|Add1~1_combout ),
	.src_payload6(\cmd_mux|src_payload~9_combout ),
	.Add31(\hps_0_h2f_lw_axi_master_agent|Add3~1_combout ),
	.src_data_71(\cmd_mux|src_data[71]~5_combout ),
	.src_payload7(\cmd_mux|src_payload~10_combout ),
	.LessThan12(\hps_0_h2f_lw_axi_master_agent|LessThan12~0_combout ),
	.src_payload8(\cmd_mux|src_payload~11_combout ),
	.src_data_72(\cmd_mux|src_data[72]~8_combout ),
	.address_burst_2(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[2]~q ),
	.src_data_38(\cmd_mux|src_data[38]~combout ),
	.src_payload9(\cmd_mux|src_payload~12_combout ),
	.src_data_73(\cmd_mux|src_data[73]~11_combout ),
	.address_burst_3(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[3]~q ),
	.src_data_39(\cmd_mux|src_data[39]~combout ),
	.src_payload10(\cmd_mux|src_payload~13_combout ),
	.src_payload11(\cmd_mux|src_payload~14_combout ),
	.src_data_74(\cmd_mux|src_data[74]~13_combout ),
	.src_payload12(\cmd_mux|src_payload~15_combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.src_data_701(\cmd_mux|src_data[70]~15_combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.src_data_711(\cmd_mux|src_data[71]~17_combout ),
	.src_data_721(\cmd_mux|src_data[72]~19_combout ),
	.src_data_731(\cmd_mux|src_data[73]~21_combout ),
	.src_payload13(\cmd_mux|src_payload~17_combout ),
	.src_data_741(\cmd_mux|src_data[74]~23_combout ),
	.clk_clk(clk_clk));

system_altera_merlin_burst_adapter ram_s1_burst_adapter(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_1(int_nxt_addr_reg_dly_1),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.out_uncomp_byte_cnt_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[1]~q ),
	.out_uncomp_byte_cnt_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[0]~q ),
	.out_uncomp_byte_cnt_reg_5(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_4(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_burstwrap_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ),
	.out_addr_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ),
	.out_burstwrap_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ),
	.out_data_49(\ram_s1_cmd_width_adapter|out_data[49]~36_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.stateST_COMP_TRANS(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.nxt_out_eop(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.in_data_reg_59(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.in_narrow_reg(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\ram_s1_agent|WideOr0~combout ),
	.in_ready_hold(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.nxt_out_eop1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.nxt_in_ready(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready2(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.in_data_reg_41(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[41]~q ),
	.source0_data_16(source0_data_16),
	.source0_data_17(source0_data_17),
	.write_addr_data_both_valid(\hps_0_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ),
	.r_sync_rst(r_sync_rst),
	.use_reg(\ram_s1_cmd_width_adapter|use_reg~q ),
	.out_endofpacket(\ram_s1_cmd_width_adapter|out_endofpacket~1_combout ),
	.out_data_59(\ram_s1_cmd_width_adapter|out_data[59]~0_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_data_70(\cmd_mux|src_data[70]~3_combout ),
	.out_data_18(\ram_s1_cmd_width_adapter|out_data[18]~2_combout ),
	.int_output_sel_0(\ram_s1_cmd_width_adapter|int_output_sel[0]~1_combout ),
	.out_data_17(\ram_s1_cmd_width_adapter|out_data[17]~3_combout ),
	.out_data_16(\ram_s1_cmd_width_adapter|out_data[16]~4_combout ),
	.in_data_reg_42(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[42]~q ),
	.out_data_50(\ram_s1_cmd_width_adapter|out_data[50]~8_combout ),
	.out_data_48(\ram_s1_cmd_width_adapter|out_data[48]~9_combout ),
	.ShiftLeft0(\ram_s1_cmd_width_adapter|ShiftLeft0~1_combout ),
	.out_data_47(\ram_s1_cmd_width_adapter|out_data[47]~10_combout ),
	.out_data_471(\ram_s1_cmd_width_adapter|out_data[47]~12_combout ),
	.out_data_51(\ram_s1_cmd_width_adapter|out_data[51]~13_combout ),
	.out_data_511(\ram_s1_cmd_width_adapter|out_data[51]~15_combout ),
	.byte_cnt_reg_1(\ram_s1_cmd_width_adapter|byte_cnt_reg[1]~q ),
	.out_data_46(\ram_s1_cmd_width_adapter|out_data[46]~16_combout ),
	.out_data_461(\ram_s1_cmd_width_adapter|out_data[46]~17_combout ),
	.cp_ready(\ram_s1_agent|cp_ready~0_combout ),
	.out_byte_cnt_reg_1(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[1]~q ),
	.in_data_reg_91(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_70(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[70]~q ),
	.in_data_reg_71(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[71]~q ),
	.in_data_reg_72(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[72]~q ),
	.in_data_reg_73(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[73]~q ),
	.in_data_reg_74(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[74]~q ),
	.in_data_reg_75(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[75]~q ),
	.in_data_reg_76(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[76]~q ),
	.in_data_reg_77(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[77]~q ),
	.in_data_reg_78(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[78]~q ),
	.in_data_reg_79(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[79]~q ),
	.in_data_reg_80(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[80]~q ),
	.in_data_reg_81(\ram_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[81]~q ),
	.out_data_0(\ram_s1_cmd_width_adapter|out_data[0]~18_combout ),
	.src_payload1(\cmd_mux|src_payload~8_combout ),
	.src_data_71(\cmd_mux|src_data[71]~5_combout ),
	.src_payload2(\cmd_mux|src_payload~10_combout ),
	.src_data_72(\cmd_mux|src_data[72]~8_combout ),
	.address_reg_2(\ram_s1_cmd_width_adapter|address_reg[2]~q ),
	.src_data_38(\cmd_mux|src_data[38]~combout ),
	.src_payload3(\cmd_mux|src_payload~12_combout ),
	.src_data_73(\cmd_mux|src_data[73]~11_combout ),
	.address_reg_3(\ram_s1_cmd_width_adapter|address_reg[3]~q ),
	.src_data_39(\cmd_mux|src_data[39]~combout ),
	.src_payload4(\cmd_mux|src_payload~13_combout ),
	.src_data_74(\cmd_mux|src_data[74]~13_combout ),
	.address_reg_4(\ram_s1_cmd_width_adapter|address_reg[4]~q ),
	.src_payload5(\cmd_mux|src_payload~15_combout ),
	.out_data_4(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~0_combout ),
	.out_data_1(\ram_s1_cmd_width_adapter|out_data[1]~19_combout ),
	.out_data_2(\ram_s1_cmd_width_adapter|out_data[2]~20_combout ),
	.out_data_3(\ram_s1_cmd_width_adapter|out_data[3]~21_combout ),
	.out_data_41(\ram_s1_cmd_width_adapter|out_data[4]~22_combout ),
	.out_data_5(\ram_s1_cmd_width_adapter|out_data[5]~23_combout ),
	.out_data_6(\ram_s1_cmd_width_adapter|out_data[6]~24_combout ),
	.out_data_7(\ram_s1_cmd_width_adapter|out_data[7]~25_combout ),
	.out_data_8(\ram_s1_cmd_width_adapter|out_data[8]~26_combout ),
	.out_data_9(\ram_s1_cmd_width_adapter|out_data[9]~27_combout ),
	.out_data_10(\ram_s1_cmd_width_adapter|out_data[10]~28_combout ),
	.out_data_11(\ram_s1_cmd_width_adapter|out_data[11]~29_combout ),
	.out_data_12(\ram_s1_cmd_width_adapter|out_data[12]~30_combout ),
	.out_data_13(\ram_s1_cmd_width_adapter|out_data[13]~31_combout ),
	.out_data_14(\ram_s1_cmd_width_adapter|out_data[14]~32_combout ),
	.out_data_15(\ram_s1_cmd_width_adapter|out_data[15]~33_combout ),
	.src_data_701(\cmd_mux|src_data[70]~15_combout ),
	.out_data_481(\ram_s1_cmd_width_adapter|out_data[48]~34_combout ),
	.out_data_512(\ram_s1_cmd_width_adapter|out_data[51]~35_combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.src_data_711(\cmd_mux|src_data[71]~17_combout ),
	.src_data_721(\cmd_mux|src_data[72]~19_combout ),
	.src_data_731(\cmd_mux|src_data[73]~21_combout ),
	.src_data_741(\cmd_mux|src_data[74]~23_combout ),
	.cp_ready1(\ram_s1_agent|cp_ready~1_combout ),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

endmodule

module system_altera_avalon_sc_fifo (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_94_0,
	mem_used_01,
	src0_valid,
	mem_0_0,
	mem_1_0,
	mem_2_0,
	mem_3_0,
	mem_4_0,
	mem_5_0,
	mem_6_0,
	mem_7_0,
	mem_8_0,
	mem_9_0,
	mem_10_0,
	mem_11_0,
	mem_12_0,
	mem_13_0,
	mem_14_0,
	mem_15_0,
	reset,
	p1_ready,
	out_valid,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_94_0;
input 	mem_used_01;
input 	src0_valid;
output 	mem_0_0;
output 	mem_1_0;
output 	mem_2_0;
output 	mem_3_0;
output 	mem_4_0;
output 	mem_5_0;
output 	mem_6_0;
output 	mem_7_0;
output 	mem_8_0;
output 	mem_9_0;
output 	mem_10_0;
output 	mem_11_0;
output 	mem_12_0;
output 	mem_13_0;
output 	mem_14_0;
output 	mem_15_0;
input 	reset;
input 	p1_ready;
input 	out_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_94_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h888F888F888F888F;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!out_valid),
	.datad(!src0_valid),
	.datae(!\read~0_combout ),
	.dataf(!\mem_used[1]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'h0C0AFFFF00000000;
defparam \mem_used[1]~2 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!out_valid),
	.datad(!p1_ready),
	.datae(!\mem_used[1]~q ),
	.dataf(!\read~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h1711F3FF77773333;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!q_a_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_used_0),
	.datad(!out_valid),
	.datae(!src0_valid),
	.dataf(!\read~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFFF3FFF5F0F0F0F0;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!q_a_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!q_a_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!q_a_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!q_a_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!q_a_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!q_a_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!q_a_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!q_a_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!q_a_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!q_a_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!q_a_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!q_a_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!q_a_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!q_a_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!q_a_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

endmodule

module system_altera_avalon_sc_fifo_1 (
	int_nxt_addr_reg_dly_1,
	out_uncomp_byte_cnt_reg_1,
	out_uncomp_byte_cnt_reg_0,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0,
	nxt_out_eop,
	in_data_reg_59,
	WideOr0,
	mem_used_1,
	nxt_out_eop1,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_94_0,
	mem_used_0,
	mem_95_0,
	comb,
	mem_39_0,
	mem_51_0,
	mem_50_0,
	mem_49_0,
	mem_48_0,
	mem_47_0,
	mem_46_0,
	mem_45_0,
	last_packet_beat,
	mem_19_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_59_0,
	mem_41_0,
	mem_70_0,
	mem_71_0,
	mem_72_0,
	mem_73_0,
	mem_74_0,
	mem_75_0,
	mem_76_0,
	mem_77_0,
	mem_78_0,
	mem_79_0,
	mem_80_0,
	mem_81_0,
	in_data_reg_41,
	m0_write,
	reset,
	p1_ready,
	sink_ready,
	in_data_reg_42,
	out_byte_cnt_reg_1,
	out_valid,
	mem_53_0,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_70,
	in_data_reg_71,
	in_data_reg_72,
	in_data_reg_73,
	in_data_reg_74,
	in_data_reg_75,
	in_data_reg_76,
	in_data_reg_77,
	in_data_reg_78,
	in_data_reg_79,
	in_data_reg_80,
	in_data_reg_81,
	mem_18_0,
	mem_52_0,
	cp_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	int_nxt_addr_reg_dly_1;
input 	out_uncomp_byte_cnt_reg_1;
input 	out_uncomp_byte_cnt_reg_0;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_burstwrap_reg_1;
input 	out_addr_reg_0;
input 	out_burstwrap_reg_0;
input 	nxt_out_eop;
input 	in_data_reg_59;
input 	WideOr0;
output 	mem_used_1;
input 	nxt_out_eop1;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_94_0;
output 	mem_used_0;
output 	mem_95_0;
input 	comb;
output 	mem_39_0;
output 	mem_51_0;
output 	mem_50_0;
output 	mem_49_0;
output 	mem_48_0;
output 	mem_47_0;
output 	mem_46_0;
output 	mem_45_0;
input 	last_packet_beat;
output 	mem_19_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_59_0;
output 	mem_41_0;
output 	mem_70_0;
output 	mem_71_0;
output 	mem_72_0;
output 	mem_73_0;
output 	mem_74_0;
output 	mem_75_0;
output 	mem_76_0;
output 	mem_77_0;
output 	mem_78_0;
output 	mem_79_0;
output 	mem_80_0;
output 	mem_81_0;
input 	in_data_reg_41;
input 	m0_write;
input 	reset;
input 	p1_ready;
input 	sink_ready;
input 	in_data_reg_42;
input 	out_byte_cnt_reg_1;
input 	out_valid;
output 	mem_53_0;
input 	in_data_reg_91;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_70;
input 	in_data_reg_71;
input 	in_data_reg_72;
input 	in_data_reg_73;
input 	in_data_reg_74;
input 	in_data_reg_75;
input 	in_data_reg_76;
input 	in_data_reg_77;
input 	in_data_reg_78;
input 	in_data_reg_79;
input 	in_data_reg_80;
input 	in_data_reg_81;
output 	mem_18_0;
output 	mem_52_0;
input 	cp_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][94]~q ;
wire \mem~0_combout ;
wire \mem~31_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][95]~q ;
wire \mem~1_combout ;
wire \mem[1][42]~q ;
wire \mem~2_combout ;
wire \mem[1][51]~q ;
wire \mem~3_combout ;
wire \mem[1][50]~q ;
wire \mem~4_combout ;
wire \mem[1][49]~q ;
wire \mem~5_combout ;
wire \mem[1][48]~q ;
wire \mem~6_combout ;
wire \mem[1][47]~q ;
wire \mem~7_combout ;
wire \mem[1][46]~q ;
wire \mem~8_combout ;
wire \mem[1][45]~q ;
wire \mem~9_combout ;
wire \mem[1][19]~q ;
wire \mem~10_combout ;
wire \mem[1][91]~q ;
wire \mem~11_combout ;
wire \mem[1][92]~q ;
wire \mem~12_combout ;
wire \mem[1][93]~q ;
wire \mem~13_combout ;
wire \mem[1][59]~q ;
wire \mem~14_combout ;
wire \mem[1][41]~q ;
wire \mem~15_combout ;
wire \mem[1][70]~q ;
wire \mem~16_combout ;
wire \mem[1][71]~q ;
wire \mem~17_combout ;
wire \mem[1][72]~q ;
wire \mem~18_combout ;
wire \mem[1][73]~q ;
wire \mem~19_combout ;
wire \mem[1][74]~q ;
wire \mem~20_combout ;
wire \mem[1][75]~q ;
wire \mem~21_combout ;
wire \mem[1][76]~q ;
wire \mem~22_combout ;
wire \mem[1][77]~q ;
wire \mem~23_combout ;
wire \mem[1][78]~q ;
wire \mem~24_combout ;
wire \mem[1][79]~q ;
wire \mem~25_combout ;
wire \mem[1][80]~q ;
wire \mem~26_combout ;
wire \mem[1][81]~q ;
wire \mem~27_combout ;
wire \mem[1][53]~q ;
wire \mem~28_combout ;
wire \mem[1][18]~q ;
wire \mem~29_combout ;
wire \mem[1][52]~q ;
wire \mem~30_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][39] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_39_0),
	.prn(vcc));
defparam \mem[0][39] .is_wysiwyg = "true";
defparam \mem[0][39] .power_up = "low";

dffeas \mem[0][51] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_51_0),
	.prn(vcc));
defparam \mem[0][51] .is_wysiwyg = "true";
defparam \mem[0][51] .power_up = "low";

dffeas \mem[0][50] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_50_0),
	.prn(vcc));
defparam \mem[0][50] .is_wysiwyg = "true";
defparam \mem[0][50] .power_up = "low";

dffeas \mem[0][49] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_49_0),
	.prn(vcc));
defparam \mem[0][49] .is_wysiwyg = "true";
defparam \mem[0][49] .power_up = "low";

dffeas \mem[0][48] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_48_0),
	.prn(vcc));
defparam \mem[0][48] .is_wysiwyg = "true";
defparam \mem[0][48] .power_up = "low";

dffeas \mem[0][47] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_47_0),
	.prn(vcc));
defparam \mem[0][47] .is_wysiwyg = "true";
defparam \mem[0][47] .power_up = "low";

dffeas \mem[0][46] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_46_0),
	.prn(vcc));
defparam \mem[0][46] .is_wysiwyg = "true";
defparam \mem[0][46] .power_up = "low";

dffeas \mem[0][45] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_45_0),
	.prn(vcc));
defparam \mem[0][45] .is_wysiwyg = "true";
defparam \mem[0][45] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][41] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_41_0),
	.prn(vcc));
defparam \mem[0][41] .is_wysiwyg = "true";
defparam \mem[0][41] .power_up = "low";

dffeas \mem[0][70] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_70_0),
	.prn(vcc));
defparam \mem[0][70] .is_wysiwyg = "true";
defparam \mem[0][70] .power_up = "low";

dffeas \mem[0][71] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_71_0),
	.prn(vcc));
defparam \mem[0][71] .is_wysiwyg = "true";
defparam \mem[0][71] .power_up = "low";

dffeas \mem[0][72] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_72_0),
	.prn(vcc));
defparam \mem[0][72] .is_wysiwyg = "true";
defparam \mem[0][72] .power_up = "low";

dffeas \mem[0][73] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_73_0),
	.prn(vcc));
defparam \mem[0][73] .is_wysiwyg = "true";
defparam \mem[0][73] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][79] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_79_0),
	.prn(vcc));
defparam \mem[0][79] .is_wysiwyg = "true";
defparam \mem[0][79] .power_up = "low";

dffeas \mem[0][80] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_80_0),
	.prn(vcc));
defparam \mem[0][80] .is_wysiwyg = "true";
defparam \mem[0][80] .power_up = "low";

dffeas \mem[0][81] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_81_0),
	.prn(vcc));
defparam \mem[0][81] .is_wysiwyg = "true";
defparam \mem[0][81] .power_up = "low";

dffeas \mem[0][53] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_53_0),
	.prn(vcc));
defparam \mem[0][53] .is_wysiwyg = "true";
defparam \mem[0][53] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][52] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_52_0),
	.prn(vcc));
defparam \mem[0][52] .is_wysiwyg = "true";
defparam \mem[0][52] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!cp_ready),
	.datab(!nxt_out_eop),
	.datac(!nxt_out_eop1),
	.datad(!in_data_reg_41),
	.datae(!m0_write),
	.dataf(!in_data_reg_42),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0000001500005555;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!sink_ready),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!WideOr0),
	.datab(!in_data_reg_42),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h1111111111111111;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem~31 (
	.dataa(!out_valid_reg),
	.datab(!in_data_reg_41),
	.datac(!\mem[1][94]~q ),
	.datad(!nxt_out_eop1),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!\mem~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "on";
defparam \mem~31 .lut_mask = 64'h05150F0F15150F0F;
defparam \mem~31 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!comb),
	.datac(!last_packet_beat),
	.datad(!out_valid),
	.datae(!p1_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBAAABABABAAABABA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!sink_ready),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3313FFFF3313FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!nxt_out_eop1),
	.datad(!\mem[1][95]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2A7F2A7F2A7F2A7F;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][42] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][42]~q ),
	.prn(vcc));
defparam \mem[1][42] .is_wysiwyg = "true";
defparam \mem[1][42] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_42),
	.datac(!\mem[1][42]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][51] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][51]~q ),
	.prn(vcc));
defparam \mem[1][51] .is_wysiwyg = "true";
defparam \mem[1][51] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][51]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][50] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][50]~q ),
	.prn(vcc));
defparam \mem[1][50] .is_wysiwyg = "true";
defparam \mem[1][50] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][50]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][49] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][49]~q ),
	.prn(vcc));
defparam \mem[1][49] .is_wysiwyg = "true";
defparam \mem[1][49] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][49]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][48] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][48]~q ),
	.prn(vcc));
defparam \mem[1][48] .is_wysiwyg = "true";
defparam \mem[1][48] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][48]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][47] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][47]~q ),
	.prn(vcc));
defparam \mem[1][47] .is_wysiwyg = "true";
defparam \mem[1][47] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!\mem[1][47]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h0257025702570257;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][46] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][46]~q ),
	.prn(vcc));
defparam \mem[1][46] .is_wysiwyg = "true";
defparam \mem[1][46] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_1),
	.datad(!out_uncomp_byte_cnt_reg_1),
	.datae(!\mem[1][46]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][45] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][45]~q ),
	.prn(vcc));
defparam \mem[1][45] .is_wysiwyg = "true";
defparam \mem[1][45] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_0),
	.datad(!\mem[1][45]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h0257025702570257;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!int_nxt_addr_reg_dly_1),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h2727272727272727;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][91]~q ),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!in_data_reg_59),
	.datab(!mem_used_1),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][41] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][41]~q ),
	.prn(vcc));
defparam \mem[1][41] .is_wysiwyg = "true";
defparam \mem[1][41] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_41),
	.datac(!\mem[1][41]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h2727272727272727;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][70] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][70]~q ),
	.prn(vcc));
defparam \mem[1][70] .is_wysiwyg = "true";
defparam \mem[1][70] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][70]~q ),
	.datac(!in_data_reg_70),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][71] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][71]~q ),
	.prn(vcc));
defparam \mem[1][71] .is_wysiwyg = "true";
defparam \mem[1][71] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][71]~q ),
	.datac(!in_data_reg_71),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][72] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][72]~q ),
	.prn(vcc));
defparam \mem[1][72] .is_wysiwyg = "true";
defparam \mem[1][72] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][72]~q ),
	.datac(!in_data_reg_72),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][73] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][73]~q ),
	.prn(vcc));
defparam \mem[1][73] .is_wysiwyg = "true";
defparam \mem[1][73] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][73]~q ),
	.datac(!in_data_reg_73),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][74]~q ),
	.datac(!in_data_reg_74),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][75]~q ),
	.datac(!in_data_reg_75),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][76]~q ),
	.datac(!in_data_reg_76),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][77]~q ),
	.datac(!in_data_reg_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][78]~q ),
	.datac(!in_data_reg_78),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][79] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][79]~q ),
	.prn(vcc));
defparam \mem[1][79] .is_wysiwyg = "true";
defparam \mem[1][79] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][79]~q ),
	.datac(!in_data_reg_79),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][80] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][80]~q ),
	.prn(vcc));
defparam \mem[1][80] .is_wysiwyg = "true";
defparam \mem[1][80] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][80]~q ),
	.datac(!in_data_reg_80),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][81] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][81]~q ),
	.prn(vcc));
defparam \mem[1][81] .is_wysiwyg = "true";
defparam \mem[1][81] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][81]~q ),
	.datac(!in_data_reg_81),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][53] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][53]~q ),
	.prn(vcc));
defparam \mem[1][53] .is_wysiwyg = "true";
defparam \mem[1][53] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][53]~q ),
	.datac(!out_burstwrap_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][18]~q ),
	.datac(!out_addr_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][52] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][52]~q ),
	.prn(vcc));
defparam \mem[1][52] .is_wysiwyg = "true";
defparam \mem[1][52] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][52]~q ),
	.datac(!out_burstwrap_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~30 .shared_arith = "off";

endmodule

module system_altera_merlin_axi_master_ni (
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	Add4,
	Add5,
	Add41,
	Add51,
	Add42,
	Add52,
	Add43,
	Add53,
	Add44,
	Add54,
	in_ready,
	nxt_out_eop,
	nxt_out_eop1,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	src_valid,
	awready,
	wready,
	write_addr_data_both_valid1,
	Add1,
	src_payload,
	Add3,
	sop_enable1,
	address_burst_0,
	address_burst_1,
	write_cp_data_69,
	burst_bytecount_5,
	Add6,
	Add2,
	burst_bytecount_4,
	Add61,
	Add21,
	burst_bytecount_3,
	Add22,
	burst_bytecount_2,
	write_cp_data_66,
	write_cp_data_67,
	write_cp_data_68,
	Add11,
	src_payload1,
	Add31,
	LessThan12,
	src_payload2,
	address_burst_2,
	address_burst_3,
	src_payload3,
	out_data_4,
	altera_reset_synchronizer_int_chain_out,
	src_payload4,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
output 	Add4;
output 	Add5;
output 	Add41;
output 	Add51;
output 	Add42;
output 	Add52;
output 	Add43;
output 	Add53;
output 	Add44;
output 	Add54;
input 	in_ready;
input 	nxt_out_eop;
input 	nxt_out_eop1;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	src_valid;
output 	awready;
output 	wready;
output 	write_addr_data_both_valid1;
output 	Add1;
input 	src_payload;
output 	Add3;
output 	sop_enable1;
output 	address_burst_0;
output 	address_burst_1;
output 	write_cp_data_69;
output 	burst_bytecount_5;
output 	Add6;
output 	Add2;
output 	burst_bytecount_4;
output 	Add61;
output 	Add21;
output 	burst_bytecount_3;
output 	Add22;
output 	burst_bytecount_2;
output 	write_cp_data_66;
output 	write_cp_data_67;
output 	write_cp_data_68;
output 	Add11;
input 	src_payload1;
output 	Add31;
output 	LessThan12;
input 	src_payload2;
output 	address_burst_2;
output 	address_burst_3;
input 	src_payload3;
output 	out_data_4;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_payload4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add4~2 ;
wire \Add5~2 ;
wire \Add4~6 ;
wire \Add5~6 ;
wire \Add4~10 ;
wire \Add5~10 ;
wire \Add4~14 ;
wire \Add5~14 ;
wire \Decoder0~0_combout ;
wire \Decoder1~0_combout ;
wire \Decoder0~1_combout ;
wire \Decoder1~1_combout ;
wire \Decoder0~2_combout ;
wire \Decoder1~2_combout ;
wire \Decoder0~3_combout ;
wire \Decoder1~3_combout ;
wire \Decoder0~4_combout ;
wire \Decoder1~4_combout ;
wire \sop_enable~0_combout ;
wire \write_cp_data[65]~4_combout ;
wire \Add7~0_combout ;
wire \burst_bytecount[6]~q ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add7~3_combout ;


system_altera_merlin_address_alignment align_address_to_size(
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.wready(wready),
	.src_payload(src_payload),
	.sop_enable(sop_enable1),
	.address_burst_0(address_burst_0),
	.address_burst_1(address_burst_1),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.address_burst_2(address_burst_2),
	.address_burst_3(address_burst_3),
	.src_payload3(src_payload3),
	.out_data_4(out_data_4),
	.Decoder0(\Decoder0~0_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Decoder01(\Decoder0~1_combout ),
	.Decoder02(\Decoder0~2_combout ),
	.Decoder03(\Decoder0~3_combout ),
	.src_payload4(src_payload4),
	.Decoder04(\Decoder0~4_combout ),
	.clk(clk_clk));

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add4),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add5),
	.cout(\Add5~2 ),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add41),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add51),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add42),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add52),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add43),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add53),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add44),
	.cout(),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h00000000000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add54),
	.cout(),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h00000000000000FF;
defparam \Add5~17 .shared_arith = "off";

cyclonev_lcell_comb \awready~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!in_ready),
	.datac(!nxt_in_ready2),
	.datad(!nxt_in_ready1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(awready),
	.sumout(),
	.cout(),
	.shareout());
defparam \awready~0 .extended_lut = "off";
defparam \awready~0 .lut_mask = 64'h0000440400004404;
defparam \awready~0 .shared_arith = "off";

cyclonev_lcell_comb \wready~0 (
	.dataa(!in_ready),
	.datab(!nxt_out_eop),
	.datac(!nxt_out_eop1),
	.datad(!nxt_in_ready),
	.datae(!nxt_in_ready1),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wready),
	.sumout(),
	.cout(),
	.shareout());
defparam \wready~0 .extended_lut = "off";
defparam \wready~0 .lut_mask = 64'h00000000AAAA002A;
defparam \wready~0 .shared_arith = "off";

cyclonev_lcell_comb write_addr_data_both_valid(
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_addr_data_both_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam write_addr_data_both_valid.extended_lut = "off";
defparam write_addr_data_both_valid.lut_mask = 64'h1111111111111111;
defparam write_addr_data_both_valid.shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(!h2f_lw_AWSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00000F003F007F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00000F003F007F00;
defparam \Add3~0 .shared_arith = "off";

dffeas sop_enable(
	.clk(clk_clk),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

cyclonev_lcell_comb \write_cp_data[69]~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!sop_enable1),
	.dataf(!\burst_bytecount[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[69]~0 .extended_lut = "off";
defparam \write_cp_data[69]~0 .lut_mask = 64'h000100000001FFFF;
defparam \write_cp_data[69]~0 .shared_arith = "off";

dffeas \burst_bytecount[5] (
	.clk(clk_clk),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

cyclonev_lcell_comb \Add6~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add6~0 .extended_lut = "off";
defparam \Add6~0 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add6~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add2~0 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(clk_clk),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

cyclonev_lcell_comb \Add6~1 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add61),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \Add6~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \Add2~1 .shared_arith = "off";

dffeas \burst_bytecount[3] (
	.clk(clk_clk),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_3),
	.prn(vcc));
defparam \burst_bytecount[3] .is_wysiwyg = "true";
defparam \burst_bytecount[3] .power_up = "low";

cyclonev_lcell_comb \Add2~2 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~2 .extended_lut = "off";
defparam \Add2~2 .lut_mask = 64'h6666666666666666;
defparam \Add2~2 .shared_arith = "off";

dffeas \burst_bytecount[2] (
	.clk(clk_clk),
	.d(\write_cp_data[65]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_2),
	.prn(vcc));
defparam \burst_bytecount[2] .is_wysiwyg = "true";
defparam \burst_bytecount[2] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[66]~1 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[66]~1 .extended_lut = "off";
defparam \write_cp_data[66]~1 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[66]~1 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[67]~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[67]~2 .extended_lut = "off";
defparam \write_cp_data[67]~2 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[67]~2 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[68]~3 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!sop_enable1),
	.dataf(!burst_bytecount_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[68]~3 .extended_lut = "off";
defparam \write_cp_data[68]~3 .lut_mask = 64'h01FE000001FEFFFF;
defparam \write_cp_data[68]~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(!h2f_lw_AWSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h3F007000C0FF8FFF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h3F007000C0FF8FFF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan12~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(!h2f_lw_AWSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan12),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan12~0 .extended_lut = "off";
defparam \LessThan12~0 .lut_mask = 64'h0F003000400080FF;
defparam \LessThan12~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h0808080808080808;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[65]~4 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_cp_data[65]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[65]~4 .extended_lut = "off";
defparam \write_cp_data[65]~4 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[65]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!\write_cp_data[65]~4_combout ),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_68),
	.datad(!write_cp_data_67),
	.datae(!write_cp_data_69),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h4000BFFF4000BFFF;
defparam \Add7~0 .shared_arith = "off";

dffeas \burst_bytecount[6] (
	.clk(clk_clk),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\burst_bytecount[6]~q ),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!\write_cp_data[65]~4_combout ),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_68),
	.datad(!write_cp_data_67),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h4B0F4B0F4B0F4B0F;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!\write_cp_data[65]~4_combout ),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_67),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h4B4B4B4B4B4B4B4B;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!\write_cp_data[65]~4_combout ),
	.datab(!write_cp_data_66),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h6666666666666666;
defparam \Add7~3 .shared_arith = "off";

endmodule

module system_altera_merlin_address_alignment (
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	wready,
	src_payload,
	sop_enable,
	address_burst_0,
	address_burst_1,
	src_payload1,
	src_payload2,
	address_burst_2,
	address_burst_3,
	src_payload3,
	out_data_4,
	Decoder0,
	reset,
	Decoder01,
	Decoder02,
	Decoder03,
	src_payload4,
	Decoder04,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	wready;
input 	src_payload;
input 	sop_enable;
output 	address_burst_0;
output 	address_burst_1;
input 	src_payload1;
input 	src_payload2;
output 	address_burst_2;
output 	address_burst_3;
input 	src_payload3;
output 	out_data_4;
input 	Decoder0;
input 	reset;
input 	Decoder01;
input 	Decoder02;
input 	Decoder03;
input 	src_payload4;
input 	Decoder04;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_data[0]~1_combout ;
wire \Add1~1_sumout ;
wire \Add0~1_sumout ;
wire \Selector20~0_combout ;
wire \out_data[1]~2_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Selector19~0_combout ;
wire \out_data[2]~3_combout ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Selector18~0_combout ;
wire \out_data[3]~4_combout ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Selector17~0_combout ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Selector16~0_combout ;
wire \address_burst[4]~q ;


dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_0),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_1),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_2),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_3),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

cyclonev_lcell_comb \out_data[4]~0 (
	.dataa(!h2f_lw_AWADDR_4),
	.datab(!sop_enable),
	.datac(!\address_burst[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~0 .extended_lut = "off";
defparam \out_data[4]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~1 (
	.dataa(!h2f_lw_AWADDR_0),
	.datab(!sop_enable),
	.datac(!address_burst_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~1 .extended_lut = "off";
defparam \out_data[0]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_0),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(!address_burst_0),
	.datac(!h2f_lw_AWADDR_0),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!Decoder0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload),
	.datad(!\out_data[0]~1_combout ),
	.datae(!\Add1~1_sumout ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector20~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~2 (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!sop_enable),
	.datac(!address_burst_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~2 .extended_lut = "off";
defparam \out_data[1]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_1),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_1),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\out_data[1]~2_combout ),
	.datad(!src_payload1),
	.datae(!\Add1~5_sumout ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector19~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[2]~3 (
	.dataa(!h2f_lw_AWADDR_2),
	.datab(!sop_enable),
	.datac(!address_burst_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~3 .extended_lut = "off";
defparam \out_data[2]~3 .lut_mask = 64'h4747474747474747;
defparam \out_data[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!address_burst_2),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!address_burst_2),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload2),
	.datad(!\out_data[2]~3_combout ),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector18~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~4 (
	.dataa(!h2f_lw_AWADDR_3),
	.datab(!sop_enable),
	.datac(!address_burst_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~4 .extended_lut = "off";
defparam \out_data[3]~4 .lut_mask = 64'h4747474747474747;
defparam \out_data[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!address_burst_3),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!address_burst_3),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload4),
	.datad(!\out_data[3]~4_combout ),
	.datae(!\Add1~13_sumout ),
	.dataf(!\Add0~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload3),
	.datad(!out_data_4),
	.datae(!\Add1~17_sumout ),
	.dataf(!\Add0~17_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector16~0 .shared_arith = "off";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[4]~q ),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

endmodule

module system_altera_merlin_burst_adapter (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	in_data_reg_0,
	int_nxt_addr_reg_dly_1,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	out_uncomp_byte_cnt_reg_1,
	out_uncomp_byte_cnt_reg_0,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0,
	out_data_49,
	saved_grant_1,
	saved_grant_0,
	src_data_78,
	src_data_79,
	src_data_77,
	stateST_COMP_TRANS,
	nxt_out_eop,
	in_data_reg_59,
	in_narrow_reg,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	in_ready_hold,
	mem_used_1,
	nxt_out_eop1,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	nxt_in_ready2,
	in_data_reg_41,
	source0_data_16,
	source0_data_17,
	write_addr_data_both_valid,
	r_sync_rst,
	use_reg,
	out_endofpacket,
	out_data_59,
	src_payload,
	src_data_70,
	out_data_18,
	int_output_sel_0,
	out_data_17,
	out_data_16,
	in_data_reg_42,
	out_data_50,
	out_data_48,
	ShiftLeft0,
	out_data_47,
	out_data_471,
	out_data_51,
	out_data_511,
	byte_cnt_reg_1,
	out_data_46,
	out_data_461,
	cp_ready,
	out_byte_cnt_reg_1,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_70,
	in_data_reg_71,
	in_data_reg_72,
	in_data_reg_73,
	in_data_reg_74,
	in_data_reg_75,
	in_data_reg_76,
	in_data_reg_77,
	in_data_reg_78,
	in_data_reg_79,
	in_data_reg_80,
	in_data_reg_81,
	out_data_0,
	src_payload1,
	src_data_71,
	src_payload2,
	src_data_72,
	address_reg_2,
	src_data_38,
	src_payload3,
	src_data_73,
	address_reg_3,
	src_data_39,
	src_payload4,
	src_data_74,
	address_reg_4,
	src_payload5,
	out_data_4,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_41,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	src_data_701,
	out_data_481,
	out_data_512,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_711,
	src_data_721,
	src_data_731,
	src_data_741,
	cp_ready1,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_1;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	out_uncomp_byte_cnt_reg_1;
output 	out_uncomp_byte_cnt_reg_0;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_burstwrap_reg_1;
output 	out_addr_reg_0;
output 	out_burstwrap_reg_0;
input 	out_data_49;
input 	saved_grant_1;
input 	saved_grant_0;
input 	src_data_78;
input 	src_data_79;
input 	src_data_77;
output 	stateST_COMP_TRANS;
output 	nxt_out_eop;
output 	in_data_reg_59;
output 	in_narrow_reg;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
output 	in_ready_hold;
input 	mem_used_1;
output 	nxt_out_eop1;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
output 	nxt_in_ready2;
output 	in_data_reg_41;
output 	source0_data_16;
output 	source0_data_17;
input 	write_addr_data_both_valid;
input 	r_sync_rst;
input 	use_reg;
input 	out_endofpacket;
input 	out_data_59;
input 	src_payload;
input 	src_data_70;
input 	out_data_18;
input 	int_output_sel_0;
input 	out_data_17;
input 	out_data_16;
output 	in_data_reg_42;
input 	out_data_50;
input 	out_data_48;
input 	ShiftLeft0;
input 	out_data_47;
input 	out_data_471;
input 	out_data_51;
input 	out_data_511;
input 	byte_cnt_reg_1;
input 	out_data_46;
input 	out_data_461;
input 	cp_ready;
output 	out_byte_cnt_reg_1;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_70;
output 	in_data_reg_71;
output 	in_data_reg_72;
output 	in_data_reg_73;
output 	in_data_reg_74;
output 	in_data_reg_75;
output 	in_data_reg_76;
output 	in_data_reg_77;
output 	in_data_reg_78;
output 	in_data_reg_79;
output 	in_data_reg_80;
output 	in_data_reg_81;
input 	out_data_0;
input 	src_payload1;
input 	src_data_71;
input 	src_payload2;
input 	src_data_72;
input 	address_reg_2;
input 	src_data_38;
input 	src_payload3;
input 	src_data_73;
input 	address_reg_3;
input 	src_data_39;
input 	src_payload4;
input 	src_data_74;
input 	address_reg_4;
input 	src_payload5;
input 	out_data_4;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_41;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	out_data_8;
input 	out_data_9;
input 	out_data_10;
input 	out_data_11;
input 	out_data_12;
input 	out_data_13;
input 	out_data_14;
input 	out_data_15;
input 	src_data_701;
input 	out_data_481;
input 	out_data_512;
input 	src_data_88;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_711;
input 	src_data_721;
input 	src_data_731;
input 	src_data_741;
input 	cp_ready1;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altera_merlin_burst_adapter_13_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_1(int_nxt_addr_reg_dly_1),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.out_uncomp_byte_cnt_reg_1(out_uncomp_byte_cnt_reg_1),
	.out_uncomp_byte_cnt_reg_0(out_uncomp_byte_cnt_reg_0),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_burstwrap_reg_1(out_burstwrap_reg_1),
	.out_addr_reg_0(out_addr_reg_0),
	.out_burstwrap_reg_0(out_burstwrap_reg_0),
	.out_data_49(out_data_49),
	.sink0_data({src_data_79,src_data_78,src_data_77,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,src_data_91,src_data_90,src_data_89,src_data_88,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_59,gnd,gnd,src_data_741,
src_data_731,src_data_721,src_data_711,src_data_701,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,
out_data_10,out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_41,out_data_3,out_data_2,out_data_1,out_data_0}),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.nxt_out_eop(nxt_out_eop),
	.in_data_reg_59(in_data_reg_59),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.WideOr0(WideOr0),
	.in_ready_hold1(in_ready_hold),
	.mem_used_1(mem_used_1),
	.nxt_out_eop1(nxt_out_eop1),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.nxt_in_ready2(nxt_in_ready2),
	.in_data_reg_41(in_data_reg_41),
	.source0_data_16(source0_data_16),
	.source0_data_17(source0_data_17),
	.write_addr_data_both_valid(write_addr_data_both_valid),
	.r_sync_rst(r_sync_rst),
	.use_reg(use_reg),
	.sink0_endofpacket(out_endofpacket),
	.src_payload(src_payload),
	.src_data_70(src_data_70),
	.out_data_18(out_data_18),
	.int_output_sel_0(int_output_sel_0),
	.in_data_reg_42(in_data_reg_42),
	.out_data_50(out_data_50),
	.out_data_48(out_data_48),
	.ShiftLeft0(ShiftLeft0),
	.out_data_47(out_data_47),
	.out_data_471(out_data_471),
	.out_data_51(out_data_51),
	.out_data_511(out_data_511),
	.byte_cnt_reg_1(byte_cnt_reg_1),
	.out_data_46(out_data_46),
	.out_data_461(out_data_461),
	.cp_ready(cp_ready),
	.out_byte_cnt_reg_1(out_byte_cnt_reg_1),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_70(in_data_reg_70),
	.in_data_reg_71(in_data_reg_71),
	.in_data_reg_72(in_data_reg_72),
	.in_data_reg_73(in_data_reg_73),
	.in_data_reg_74(in_data_reg_74),
	.in_data_reg_75(in_data_reg_75),
	.in_data_reg_76(in_data_reg_76),
	.in_data_reg_77(in_data_reg_77),
	.in_data_reg_78(in_data_reg_78),
	.in_data_reg_79(in_data_reg_79),
	.in_data_reg_80(in_data_reg_80),
	.in_data_reg_81(in_data_reg_81),
	.src_payload1(src_payload1),
	.src_data_71(src_data_71),
	.src_payload2(src_payload2),
	.src_data_72(src_data_72),
	.address_reg_2(address_reg_2),
	.src_data_38(src_data_38),
	.src_payload3(src_payload3),
	.src_data_73(src_data_73),
	.address_reg_3(address_reg_3),
	.src_data_39(src_data_39),
	.src_payload4(src_payload4),
	.src_data_74(src_data_74),
	.address_reg_4(address_reg_4),
	.src_payload5(src_payload5),
	.out_data_4(out_data_4),
	.out_data_481(out_data_481),
	.out_data_512(out_data_512),
	.cp_ready1(cp_ready1),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

endmodule

module system_altera_merlin_burst_adapter_13_1 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	in_data_reg_0,
	int_nxt_addr_reg_dly_1,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	out_uncomp_byte_cnt_reg_1,
	out_uncomp_byte_cnt_reg_0,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0,
	out_data_49,
	sink0_data,
	stateST_COMP_TRANS,
	nxt_out_eop,
	in_data_reg_59,
	in_narrow_reg1,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	in_ready_hold1,
	mem_used_1,
	nxt_out_eop1,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	nxt_in_ready2,
	in_data_reg_41,
	source0_data_16,
	source0_data_17,
	write_addr_data_both_valid,
	r_sync_rst,
	use_reg,
	sink0_endofpacket,
	src_payload,
	src_data_70,
	out_data_18,
	int_output_sel_0,
	in_data_reg_42,
	out_data_50,
	out_data_48,
	ShiftLeft0,
	out_data_47,
	out_data_471,
	out_data_51,
	out_data_511,
	byte_cnt_reg_1,
	out_data_46,
	out_data_461,
	cp_ready,
	out_byte_cnt_reg_1,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_70,
	in_data_reg_71,
	in_data_reg_72,
	in_data_reg_73,
	in_data_reg_74,
	in_data_reg_75,
	in_data_reg_76,
	in_data_reg_77,
	in_data_reg_78,
	in_data_reg_79,
	in_data_reg_80,
	in_data_reg_81,
	src_payload1,
	src_data_71,
	src_payload2,
	src_data_72,
	address_reg_2,
	src_data_38,
	src_payload3,
	src_data_73,
	address_reg_3,
	src_data_39,
	src_payload4,
	src_data_74,
	address_reg_4,
	src_payload5,
	out_data_4,
	out_data_481,
	out_data_512,
	cp_ready1,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_1;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	out_uncomp_byte_cnt_reg_1;
output 	out_uncomp_byte_cnt_reg_0;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_burstwrap_reg_1;
output 	out_addr_reg_0;
output 	out_burstwrap_reg_0;
input 	out_data_49;
input 	[93:0] sink0_data;
output 	stateST_COMP_TRANS;
output 	nxt_out_eop;
output 	in_data_reg_59;
output 	in_narrow_reg1;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
output 	in_ready_hold1;
input 	mem_used_1;
output 	nxt_out_eop1;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
output 	nxt_in_ready2;
output 	in_data_reg_41;
output 	source0_data_16;
output 	source0_data_17;
input 	write_addr_data_both_valid;
input 	r_sync_rst;
input 	use_reg;
input 	sink0_endofpacket;
input 	src_payload;
input 	src_data_70;
input 	out_data_18;
input 	int_output_sel_0;
output 	in_data_reg_42;
input 	out_data_50;
input 	out_data_48;
input 	ShiftLeft0;
input 	out_data_47;
input 	out_data_471;
input 	out_data_51;
input 	out_data_511;
input 	byte_cnt_reg_1;
input 	out_data_46;
input 	out_data_461;
input 	cp_ready;
output 	out_byte_cnt_reg_1;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_70;
output 	in_data_reg_71;
output 	in_data_reg_72;
output 	in_data_reg_73;
output 	in_data_reg_74;
output 	in_data_reg_75;
output 	in_data_reg_76;
output 	in_data_reg_77;
output 	in_data_reg_78;
output 	in_data_reg_79;
output 	in_data_reg_80;
output 	in_data_reg_81;
input 	src_payload1;
input 	src_data_71;
input 	src_payload2;
input 	src_data_72;
input 	address_reg_2;
input 	src_data_38;
input 	src_payload3;
input 	src_data_73;
input 	address_reg_3;
input 	src_data_39;
input 	src_payload4;
input 	src_data_74;
input 	address_reg_4;
input 	src_payload5;
input 	out_data_4;
input 	out_data_481;
input 	out_data_512;
input 	cp_ready1;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|out_data[0]~combout ;
wire \in_valid~combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_eop_reg~q ;
wire \Add4~6 ;
wire \Add4~7 ;
wire \Add4~14 ;
wire \Add4~15 ;
wire \Add4~10 ;
wire \Add4~11 ;
wire \Add4~26 ;
wire \Add4~27 ;
wire \Add4~22 ;
wire \Add4~23 ;
wire \Add4~18 ;
wire \Add4~19 ;
wire \Add4~1_sumout ;
wire \Selector3~0_combout ;
wire \Add4~5_sumout ;
wire \Add4~9_sumout ;
wire \Add4~13_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[1]~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~5_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~6_combout ;
wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \Add4~17_sumout ;
wire \Add4~21_sumout ;
wire \Add4~25_sumout ;
wire \WideOr0~2_combout ;
wire \new_burst_reg~0_combout ;
wire \WideNor0~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_eop~2_combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \Selector2~3_combout ;
wire \Selector2~4_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \nxt_in_ready~1_combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \new_burst_reg~1_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \Add1~21_sumout ;
wire \int_bytes_remaining_reg[0]~q ;
wire \Add1~22 ;
wire \Add1~23 ;
wire \Add1~25_sumout ;
wire \int_bytes_remaining_reg[1]~q ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~1_sumout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~2 ;
wire \Add1~3 ;
wire \Add1~5_sumout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~6 ;
wire \Add1~7 ;
wire \Add1~9_sumout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~10 ;
wire \Add1~11 ;
wire \Add1~13_sumout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \Add1~14 ;
wire \Add1~15 ;
wire \Add1~17_sumout ;
wire \new_burst_reg~2_combout ;
wire \new_burst_reg~3_combout ;
wire \new_burst_reg~4_combout ;
wire \new_burst_reg~q ;
wire \d0_in_size[0]~0_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~0_combout ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \int_nxt_addr_with_offset[0]~combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~1_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \int_nxt_addr_with_offset[1]~combout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \d0_int_nxt_addr[2]~0_combout ;
wire \nxt_addr[2]~2_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \int_nxt_addr_with_offset[2]~combout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \d0_int_nxt_addr[3]~1_combout ;
wire \nxt_addr[3]~3_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \int_nxt_addr_with_offset[3]~combout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \in_burstwrap_reg[4]~q ;
wire \d0_int_nxt_addr[4]~2_combout ;
wire \nxt_addr[4]~4_combout ;
wire \int_nxt_addr_reg[4]~q ;
wire \int_nxt_addr_with_offset[4]~combout ;
wire \always10~0_combout ;
wire \in_narrow_reg~0_combout ;
wire \nxt_out_valid~0_combout ;
wire \WideOr0~5_combout ;
wire \WideOr0~3_combout ;
wire \WideOr0~4_combout ;
wire \Selector3~1_combout ;


system_altera_merlin_address_alignment_1 align_address_to_size(
	.d0_in_size_0(\d0_in_size[0]~0_combout ),
	.out_data_18(out_data_18),
	.out_data_0(\align_address_to_size|out_data[0]~combout ));

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\int_nxt_addr_with_offset[1]~combout ),
	.asdata(int_output_sel_0),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_1),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\int_nxt_addr_with_offset[2]~combout ),
	.asdata(\d0_int_nxt_addr[2]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\int_nxt_addr_with_offset[3]~combout ),
	.asdata(\d0_int_nxt_addr[3]~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[4] (
	.clk(clk_clk),
	.d(\int_nxt_addr_with_offset[4]~combout ),
	.asdata(\d0_int_nxt_addr[4]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_4),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[4] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(clk_clk),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(clk_clk),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(clk_clk),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(clk_clk),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(clk_clk),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(clk_clk),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(clk_clk),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(clk_clk),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(clk_clk),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!sink0_data[41]),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[1] (
	.clk(clk_clk),
	.d(\Add4~13_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[1]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_1),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[1] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[1] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[0] (
	.clk(clk_clk),
	.d(\Add4~5_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_0),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[0] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[0] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\Add4~17_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\Add4~1_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\Add4~21_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\Add4~25_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[3]~5_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\Add4~9_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[2]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(\in_burstwrap_reg[1]~q ),
	.asdata(sink0_data[53]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\always10~0_combout ),
	.q(out_burstwrap_reg_1),
	.prn(vcc));
defparam \out_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[1] .power_up = "low";

dffeas \out_addr_reg[0] (
	.clk(clk_clk),
	.d(\int_nxt_addr_with_offset[0]~combout ),
	.asdata(out_data_18),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_addr_reg_0),
	.prn(vcc));
defparam \out_addr_reg[0] .is_wysiwyg = "true";
defparam \out_addr_reg[0] .power_up = "low";

dffeas \out_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(\in_burstwrap_reg[0]~q ),
	.asdata(sink0_data[52]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\always10~0_combout ),
	.q(out_burstwrap_reg_0),
	.prn(vcc));
defparam \out_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[0] .power_up = "low";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\in_eop_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h2222222222222222;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[59] (
	.clk(clk_clk),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\in_narrow_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas in_ready_hold(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_hold1),
	.prn(vcc));
defparam in_ready_hold.is_wysiwyg = "true";
defparam in_ready_hold.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!\new_burst_reg~q ),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~1 .extended_lut = "off";
defparam \nxt_out_eop~1 .lut_mask = 64'h0000150040555555;
defparam \nxt_out_eop~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h1500150015001500;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!out_valid_reg1),
	.datab(!stateST_COMP_TRANS),
	.datac(!WideOr0),
	.datad(!in_ready_hold1),
	.datae(!mem_used_1),
	.dataf(!\nxt_in_ready~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h51115555DD11DD11;
defparam \nxt_in_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~3 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!mem_used_1),
	.datad(gnd),
	.datae(!\new_burst_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~3 .extended_lut = "off";
defparam \nxt_in_ready~3 .lut_mask = 64'h0000101000001010;
defparam \nxt_in_ready~3 .shared_arith = "off";

dffeas \in_data_reg[41] (
	.clk(clk_clk),
	.d(sink0_data[41]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_41),
	.prn(vcc));
defparam \in_data_reg[41] .is_wysiwyg = "true";
defparam \in_data_reg[41] .power_up = "low";

cyclonev_lcell_comb \source0_data[16]~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\int_nxt_addr_reg_dly[0]~q ),
	.datac(!in_narrow_reg1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[16]~0 .extended_lut = "off";
defparam \source0_data[16]~0 .lut_mask = 64'h04FE04FE04FE04FE;
defparam \source0_data[16]~0 .shared_arith = "off";

cyclonev_lcell_comb \source0_data[17]~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_data_reg_59),
	.datac(!\int_nxt_addr_reg_dly[0]~q ),
	.datad(!in_narrow_reg1),
	.datae(!in_byteen_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[17]~1 .extended_lut = "off";
defparam \source0_data[17]~1 .lut_mask = 64'h0015FFBF0015FFBF;
defparam \source0_data[17]~1 .shared_arith = "off";

dffeas \in_data_reg[42] (
	.clk(clk_clk),
	.d(sink0_data[42]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_42),
	.prn(vcc));
defparam \in_data_reg[42] .is_wysiwyg = "true";
defparam \in_data_reg[42] .power_up = "low";

dffeas \out_byte_cnt_reg[1] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_1),
	.prn(vcc));
defparam \out_byte_cnt_reg[1] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[1] .power_up = "low";

dffeas \in_data_reg[91] (
	.clk(clk_clk),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[70] (
	.clk(clk_clk),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_70),
	.prn(vcc));
defparam \in_data_reg[70] .is_wysiwyg = "true";
defparam \in_data_reg[70] .power_up = "low";

dffeas \in_data_reg[71] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_71),
	.prn(vcc));
defparam \in_data_reg[71] .is_wysiwyg = "true";
defparam \in_data_reg[71] .power_up = "low";

dffeas \in_data_reg[72] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_72),
	.prn(vcc));
defparam \in_data_reg[72] .is_wysiwyg = "true";
defparam \in_data_reg[72] .power_up = "low";

dffeas \in_data_reg[73] (
	.clk(clk_clk),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_73),
	.prn(vcc));
defparam \in_data_reg[73] .is_wysiwyg = "true";
defparam \in_data_reg[73] .power_up = "low";

dffeas \in_data_reg[74] (
	.clk(clk_clk),
	.d(sink0_data[74]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_74),
	.prn(vcc));
defparam \in_data_reg[74] .is_wysiwyg = "true";
defparam \in_data_reg[74] .power_up = "low";

dffeas \in_data_reg[75] (
	.clk(clk_clk),
	.d(sink0_data[75]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_75),
	.prn(vcc));
defparam \in_data_reg[75] .is_wysiwyg = "true";
defparam \in_data_reg[75] .power_up = "low";

dffeas \in_data_reg[76] (
	.clk(clk_clk),
	.d(sink0_data[76]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_76),
	.prn(vcc));
defparam \in_data_reg[76] .is_wysiwyg = "true";
defparam \in_data_reg[76] .power_up = "low";

dffeas \in_data_reg[77] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_77),
	.prn(vcc));
defparam \in_data_reg[77] .is_wysiwyg = "true";
defparam \in_data_reg[77] .power_up = "low";

dffeas \in_data_reg[78] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_78),
	.prn(vcc));
defparam \in_data_reg[78] .is_wysiwyg = "true";
defparam \in_data_reg[78] .power_up = "low";

dffeas \in_data_reg[79] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_79),
	.prn(vcc));
defparam \in_data_reg[79] .is_wysiwyg = "true";
defparam \in_data_reg[79] .power_up = "low";

dffeas \in_data_reg[80] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_80),
	.prn(vcc));
defparam \in_data_reg[80] .is_wysiwyg = "true";
defparam \in_data_reg[80] .power_up = "low";

dffeas \in_data_reg[81] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_81),
	.prn(vcc));
defparam \in_data_reg[81] .is_wysiwyg = "true";
defparam \in_data_reg[81] .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!sink0_data[42]),
	.datae(!sink0_data[41]),
	.dataf(!in_ready_hold1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000000550357;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!nxt_out_eop),
	.datab(!nxt_out_eop1),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(!\in_valid~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0000FF070000FF07;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!out_uncomp_byte_cnt_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout(\Add4~7 ));
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h0000FFFF00000F0F;
defparam \Add4~5 .shared_arith = "on";

cyclonev_lcell_comb \Add4~13 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(!out_uncomp_byte_cnt_reg_1),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(\Add4~7 ),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout(\Add4~15 ));
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000E0F0000E1F0;
defparam \Add4~13 .shared_arith = "on";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(\Add4~15 ),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout(\Add4~11 ));
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~9 .shared_arith = "on";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(\Add4~11 ),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(\Add4~26 ),
	.shareout(\Add4~27 ));
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~25 .shared_arith = "on";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~26 ),
	.sharein(\Add4~27 ),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(\Add4~22 ),
	.shareout(\Add4~23 ));
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~21 .shared_arith = "on";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(\Add4~23 ),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout(\Add4~19 ));
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~17 .shared_arith = "on";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(\Add4~19 ),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h000000000000FF00;
defparam \Add4~1 .shared_arith = "on";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!nxt_out_eop1),
	.datac(!\nxt_in_ready~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[1]~0 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_byte_cnt_reg_1),
	.dataf(!out_uncomp_byte_cnt_reg_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[1]~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[1]~0 .lut_mask = 64'h15000000FFFFEAFF;
defparam \nxt_uncomp_subburst_byte_cnt[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~1 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_uncomp_byte_cnt_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~1 .lut_mask = 64'h0000EAFF0000EAFF;
defparam \nxt_uncomp_subburst_byte_cnt~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_byte_cnt_reg_1),
	.dataf(!out_uncomp_byte_cnt_reg_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h15000000FFFFEAFF;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~3 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_byte_cnt_reg_1),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~3 .lut_mask = 64'h15000000FFFFEAFF;
defparam \nxt_uncomp_subburst_byte_cnt[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~4 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_byte_cnt_reg_1),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .lut_mask = 64'h15000000FFFFEAFF;
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~5 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_byte_cnt_reg_1),
	.dataf(!out_uncomp_byte_cnt_reg_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~5 .lut_mask = 64'h15000000FFFFEAFF;
defparam \nxt_uncomp_subburst_byte_cnt[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~6 (
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(!out_byte_cnt_reg_1),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~6 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~6 .lut_mask = 64'h15000000FFFFEAFF;
defparam \nxt_uncomp_subburst_byte_cnt[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[3]~5_combout ),
	.dataf(!\nxt_uncomp_subburst_byte_cnt[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h8000000000000000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~5_sumout ),
	.datac(!\Add4~9_sumout ),
	.datad(!\Add4~13_sumout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[1]~0_combout ),
	.dataf(!\WideOr0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'h80008000D5558000;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~17_sumout ),
	.datac(!\Add4~21_sumout ),
	.datad(!\Add4~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!out_data_48),
	.datab(!ShiftLeft0),
	.datac(!out_data_47),
	.datad(!out_data_471),
	.datae(!out_data_51),
	.dataf(!out_data_511),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hA800000000000000;
defparam \new_burst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb WideNor0(
	.dataa(!out_data_461),
	.datab(!out_data_49),
	.datac(!out_data_50),
	.datad(!\new_burst_reg~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor0.extended_lut = "off";
defparam WideNor0.lut_mask = 64'h0080008000800080;
defparam WideNor0.shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~2 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!mem_used_1),
	.datad(!\in_eop_reg~q ),
	.datae(!\new_burst_reg~q ),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_eop~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~2 .extended_lut = "off";
defparam \nxt_out_eop~2 .lut_mask = 64'h00AA10BA45EF55FF;
defparam \nxt_out_eop~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[42]),
	.datab(!sink0_data[41]),
	.datac(!nxt_out_eop),
	.datad(!nxt_out_eop1),
	.datae(!\in_valid~combout ),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h00007777F000FFFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!in_ready_hold1),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBFAABFAABFAABFAA;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!sink0_data[42]),
	.datac(!sink0_data[41]),
	.datad(!in_ready_hold1),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!write_addr_data_both_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h000000110000001F;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!sink0_data[41]),
	.datad(!in_ready_hold1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h0001000100010001;
defparam \Selector2~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~3 (
	.dataa(!sink0_data[42]),
	.datab(!\nxt_out_eop~2_combout ),
	.datac(!\state.ST_IDLE~q ),
	.datad(!\Selector2~0_combout ),
	.datae(!\Selector2~1_combout ),
	.dataf(!\Selector2~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~3 .extended_lut = "off";
defparam \Selector2~3 .lut_mask = 64'h00002222A2A0A2A2;
defparam \Selector2~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~1_sumout ),
	.datac(!\Selector3~0_combout ),
	.datad(!\WideOr0~1_combout ),
	.datae(!\WideOr0~2_combout ),
	.dataf(!\Selector2~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~4 .extended_lut = "off";
defparam \Selector2~4 .lut_mask = 64'h000D0000FFFFFFFF;
defparam \Selector2~4 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[42]),
	.datab(!sink0_data[41]),
	.datac(!stateST_COMP_TRANS),
	.datad(!\in_eop_reg~q ),
	.datae(!\nxt_in_ready~1_combout ),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hA2A2A2A2F2A2F2F2;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(gnd),
	.datac(!nxt_out_eop1),
	.datad(!\in_valid~combout ),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h50FF505050FF5050;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!use_reg),
	.datac(!byte_cnt_reg_1),
	.datad(!out_data_46),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~1 .extended_lut = "off";
defparam \new_burst_reg~1 .lut_mask = 64'h0145014501450145;
defparam \new_burst_reg~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\Add1~1_sumout ),
	.asdata(out_data_471),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout(\Add1~23 ));
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[0] (
	.clk(clk_clk),
	.d(\Add1~21_sumout ),
	.asdata(GND_port),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[0]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[0] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!out_byte_cnt_reg_1),
	.datad(!\int_bytes_remaining_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(\Add1~23 ),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout(\Add1~27 ));
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000F00000F00F;
defparam \Add1~25 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[1] (
	.clk(clk_clk),
	.d(\Add1~25_sumout ),
	.asdata(out_data_461),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[1]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[1] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[1] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(\Add1~27 ),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout(\Add1~3 ));
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~1 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\Add1~5_sumout ),
	.asdata(out_data_481),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(\Add1~3 ),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout(\Add1~7 ));
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~5 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\Add1~9_sumout ),
	.asdata(out_data_49),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(\Add1~7 ),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout(\Add1~11 ));
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~9 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\Add1~13_sumout ),
	.asdata(out_data_50),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(\Add1~11 ),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout(\Add1~15 ));
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~13 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\Add1~17_sumout ),
	.asdata(out_data_512),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(\Add1~15 ),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "on";

cyclonev_lcell_comb \new_burst_reg~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add1~21_sumout ),
	.datac(!\Add1~25_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~2 .extended_lut = "off";
defparam \new_burst_reg~2 .lut_mask = 64'h0808080808080808;
defparam \new_burst_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~3 (
	.dataa(!\Add1~1_sumout ),
	.datab(!\Add1~5_sumout ),
	.datac(!\Add1~9_sumout ),
	.datad(!\Add1~13_sumout ),
	.datae(!\Add1~17_sumout ),
	.dataf(!\new_burst_reg~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~3 .extended_lut = "off";
defparam \new_burst_reg~3 .lut_mask = 64'h0000000080000000;
defparam \new_burst_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~4 (
	.dataa(!\Selector1~1_combout ),
	.datab(!out_data_49),
	.datac(!out_data_50),
	.datad(!\new_burst_reg~0_combout ),
	.datae(!\new_burst_reg~1_combout ),
	.dataf(!\new_burst_reg~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~4 .extended_lut = "off";
defparam \new_burst_reg~4 .lut_mask = 64'hAAAAAAEAFFFFFFFF;
defparam \new_burst_reg~4 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \d0_in_size[0]~0 (
	.dataa(!sink0_data[92]),
	.datab(!sink0_data[93]),
	.datac(!sink0_data[91]),
	.datad(!in_data_reg_59),
	.datae(!\new_burst_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_in_size[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_in_size[0]~0 .extended_lut = "off";
defparam \d0_in_size[0]~0 .lut_mask = 64'h00FF7F7F00FF7F7F;
defparam \d0_in_size[0]~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\d0_in_size[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

cyclonev_lcell_comb \int_byte_cnt_narrow_reg[0]~0 (
	.dataa(!\d0_in_size[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_byte_cnt_narrow_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_byte_cnt_narrow_reg[0]~0 .extended_lut = "off";
defparam \int_byte_cnt_narrow_reg[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \int_byte_cnt_narrow_reg[0]~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\int_byte_cnt_narrow_reg[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[52]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(gnd),
	.datac(!sink0_data[52]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\align_address_to_size|out_data[0]~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "off";
defparam \nxt_addr[0]~0 .lut_mask = 64'h0000AA005050FA50;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~1_sumout ),
	.datac(!src_payload),
	.datad(!src_data_70),
	.datae(!\in_burstwrap_reg[0]~q ),
	.dataf(!\int_nxt_addr_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[0] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[0] .lut_mask = 64'h11013323FFFFFFFF;
defparam \int_nxt_addr_with_offset[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\int_nxt_addr_with_offset[0]~combout ),
	.asdata(\align_address_to_size|out_data[0]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\new_burst_reg~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_1),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[53]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!int_output_sel_0),
	.datac(gnd),
	.datad(!sink0_data[53]),
	.datae(!\in_burstwrap_reg[1]~q ),
	.dataf(!\int_nxt_addr_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~1 .extended_lut = "off";
defparam \nxt_addr[1]~1 .lut_mask = 64'h11001100BBAA1100;
defparam \nxt_addr[1]~1 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~5_sumout ),
	.datac(!src_payload1),
	.datad(!src_data_71),
	.datae(!\in_burstwrap_reg[1]~q ),
	.dataf(!\int_nxt_addr_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[1] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[1] .lut_mask = 64'h11013323FFFFFFFF;
defparam \int_nxt_addr_with_offset[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[54]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~0 (
	.dataa(!use_reg),
	.datab(!address_reg_2),
	.datac(!src_data_38),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \d0_int_nxt_addr[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(gnd),
	.datac(!sink0_data[54]),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\int_nxt_addr_reg[2]~q ),
	.dataf(!\d0_int_nxt_addr[2]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~2 .extended_lut = "off";
defparam \nxt_addr[2]~2 .lut_mask = 64'h0000AA005050FA50;
defparam \nxt_addr[2]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!src_payload2),
	.datad(!src_data_72),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\int_nxt_addr_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[2] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[2] .lut_mask = 64'h11013323FFFFFFFF;
defparam \int_nxt_addr_with_offset[2] .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[55]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~1 (
	.dataa(!use_reg),
	.datab(!address_reg_3),
	.datac(!src_data_39),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \d0_int_nxt_addr[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(gnd),
	.datac(!sink0_data[55]),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\int_nxt_addr_reg[3]~q ),
	.dataf(!\d0_int_nxt_addr[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~3 .extended_lut = "off";
defparam \nxt_addr[3]~3 .lut_mask = 64'h0000AA005050FA50;
defparam \nxt_addr[3]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!src_payload3),
	.datad(!src_data_73),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\int_nxt_addr_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[3] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[3] .lut_mask = 64'h11013323FFFFFFFF;
defparam \int_nxt_addr_with_offset[3] .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \in_burstwrap_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[56]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[4]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[4] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~2 (
	.dataa(!sink0_data[41]),
	.datab(!use_reg),
	.datac(!address_reg_4),
	.datad(!src_payload5),
	.datae(!out_data_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~2 .lut_mask = 64'h03CF47CF03CF47CF;
defparam \d0_int_nxt_addr[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[4]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(gnd),
	.datac(!sink0_data[56]),
	.datad(!\in_burstwrap_reg[4]~q ),
	.datae(!\int_nxt_addr_reg[4]~q ),
	.dataf(!\d0_int_nxt_addr[4]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[4]~4 .extended_lut = "off";
defparam \nxt_addr[4]~4 .lut_mask = 64'h0000AA005050FA50;
defparam \nxt_addr[4]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[4] (
	.clk(clk_clk),
	.d(\nxt_addr[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[4]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[4] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[4] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~17_sumout ),
	.datac(!src_payload4),
	.datad(!src_data_74),
	.datae(!\in_burstwrap_reg[4]~q ),
	.dataf(!\int_nxt_addr_reg[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[4] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[4] .lut_mask = 64'h11013323FFFFFFFF;
defparam \int_nxt_addr_with_offset[4] .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!out_valid_reg1),
	.datab(!stateST_COMP_TRANS),
	.datac(!cp_ready1),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(!nxt_out_eop1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'hAEAAAEAAAFAAAFAA;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \in_narrow_reg~0 (
	.dataa(!sink0_data[59]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_narrow_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_narrow_reg~0 .extended_lut = "off";
defparam \in_narrow_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_narrow_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~17_sumout ),
	.datac(!\Add4~1_sumout ),
	.datad(!\Add4~21_sumout ),
	.datae(!\Add4~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~5 .extended_lut = "off";
defparam \WideOr0~5 .lut_mask = 64'h2AAAAAAA2AAAAAAA;
defparam \WideOr0~5 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready1),
	.datac(!mem_used_1),
	.datad(!out_byte_cnt_reg_1),
	.datae(!out_uncomp_byte_cnt_reg_0),
	.dataf(!out_uncomp_byte_cnt_reg_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'hEFFF001000100010;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~5_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~6_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[1]~0_combout ),
	.dataf(!\WideOr0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\Add4~5_sumout ),
	.datab(!\WideOr0~5_combout ),
	.datac(!\WideOr0~4_combout ),
	.datad(!\Selector3~0_combout ),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!\Add4~9_sumout ),
	.datag(!\Add4~13_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "on";
defparam \Selector3~1 .lut_mask = 64'h007F003F00FF003F;
defparam \Selector3~1 .shared_arith = "off";

endmodule

module system_altera_merlin_address_alignment_1 (
	d0_in_size_0,
	out_data_18,
	out_data_0)/* synthesis synthesis_greybox=0 */;
input 	d0_in_size_0;
input 	out_data_18;
output 	out_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \out_data[0] (
	.dataa(!d0_in_size_0),
	.datab(!out_data_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0] .extended_lut = "off";
defparam \out_data[0] .lut_mask = 64'h2222222222222222;
defparam \out_data[0] .shared_arith = "off";

endmodule

module system_altera_merlin_slave_agent (
	always10,
	stateST_COMP_TRANS,
	in_narrow_reg,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr01,
	in_ready_hold,
	mem_used_1,
	out_valid_reg,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_94_0,
	mem_used_01,
	out_valid,
	mem_95_0,
	comb,
	mem_39_0,
	mem_51_0,
	mem_50_0,
	mem_49_0,
	mem_48_0,
	mem_47_0,
	mem_46_0,
	mem_45_0,
	last_packet_beat,
	source_addr_1,
	source_addr_11,
	mem_19_0,
	mem_59_0,
	source_endofpacket,
	in_data_reg_41,
	m0_write,
	m0_write1,
	r_sync_rst,
	p1_ready,
	rf_sink_ready,
	cp_ready,
	out_valid1,
	mem_53_0,
	mem_18_0,
	mem_52_0,
	cp_ready1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	always10;
input 	stateST_COMP_TRANS;
input 	in_narrow_reg;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr01;
input 	in_ready_hold;
input 	mem_used_1;
input 	out_valid_reg;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_94_0;
input 	mem_used_01;
input 	out_valid;
input 	mem_95_0;
output 	comb;
input 	mem_39_0;
input 	mem_51_0;
input 	mem_50_0;
input 	mem_49_0;
input 	mem_48_0;
input 	mem_47_0;
input 	mem_46_0;
input 	mem_45_0;
output 	last_packet_beat;
output 	source_addr_1;
output 	source_addr_11;
input 	mem_19_0;
input 	mem_59_0;
output 	source_endofpacket;
input 	in_data_reg_41;
output 	m0_write;
output 	m0_write1;
input 	r_sync_rst;
input 	p1_ready;
output 	rf_sink_ready;
output 	cp_ready;
input 	out_valid1;
input 	mem_53_0;
input 	mem_18_0;
input 	mem_52_0;
output 	cp_ready1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altera_merlin_burst_uncompressor uncompressor(
	.always10(always10),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_used_0(mem_used_0),
	.mem_94_0(mem_94_0),
	.mem_used_01(mem_used_01),
	.out_valid(out_valid),
	.mem_95_0(mem_95_0),
	.comb(comb),
	.mem_39_0(mem_39_0),
	.mem_51_0(mem_51_0),
	.mem_50_0(mem_50_0),
	.mem_49_0(mem_49_0),
	.mem_48_0(mem_48_0),
	.mem_47_0(mem_47_0),
	.mem_46_0(mem_46_0),
	.mem_45_0(mem_45_0),
	.last_packet_beat(last_packet_beat),
	.source_addr_1(source_addr_1),
	.source_addr_11(source_addr_11),
	.mem_19_0(mem_19_0),
	.mem_59_0(mem_59_0),
	.source_endofpacket1(source_endofpacket),
	.reset(r_sync_rst),
	.p1_ready(p1_ready),
	.sink_ready(rf_sink_ready),
	.out_valid1(out_valid1),
	.mem_53_0(mem_53_0),
	.mem_18_0(mem_18_0),
	.mem_52_0(mem_52_0),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr0(
	.dataa(!stateST_COMP_TRANS),
	.datab(gnd),
	.datac(gnd),
	.datad(!in_narrow_reg),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'hFFAA000000000000;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_94_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~0 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'h4444444444444444;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!WideOr01),
	.datab(!in_data_reg_41),
	.datac(!m0_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'h0202020202020202;
defparam \m0_write~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_narrow_reg),
	.datab(!in_byteen_reg_1),
	.datac(!in_byteen_reg_0),
	.datad(!in_ready_hold),
	.datae(!mem_used_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h80FF000080FF0000;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_narrow_reg),
	.datab(!stateST_COMP_TRANS),
	.datac(!in_ready_hold),
	.datad(!in_byteen_reg_0),
	.datae(!in_byteen_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'hEF0F0F0FEF0F0F0F;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module system_altera_merlin_burst_uncompressor (
	always10,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_94_0,
	mem_used_01,
	out_valid,
	mem_95_0,
	comb,
	mem_39_0,
	mem_51_0,
	mem_50_0,
	mem_49_0,
	mem_48_0,
	mem_47_0,
	mem_46_0,
	mem_45_0,
	last_packet_beat,
	source_addr_1,
	source_addr_11,
	mem_19_0,
	mem_59_0,
	source_endofpacket1,
	reset,
	p1_ready,
	sink_ready,
	out_valid1,
	mem_53_0,
	mem_18_0,
	mem_52_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	always10;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_94_0;
input 	mem_used_01;
input 	out_valid;
input 	mem_95_0;
input 	comb;
input 	mem_39_0;
input 	mem_51_0;
input 	mem_50_0;
input 	mem_49_0;
input 	mem_48_0;
input 	mem_47_0;
input 	mem_46_0;
input 	mem_45_0;
output 	last_packet_beat;
output 	source_addr_1;
output 	source_addr_11;
input 	mem_19_0;
input 	mem_59_0;
output 	source_endofpacket1;
input 	reset;
input 	p1_ready;
output 	sink_ready;
input 	out_valid1;
input 	mem_53_0;
input 	mem_18_0;
input 	mem_52_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \Add0~3_combout ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \Add1~2_combout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~1_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \burst_uncompress_byte_counter~7_combout ;
wire \burst_uncompress_byte_counter[0]~q ;
wire \last_packet_beat~1_combout ;
wire \burst_uncompress_byte_counter~8_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[1]~q ;
wire \last_packet_beat~0_combout ;
wire \last_packet_beat~2_combout ;
wire \last_packet_beat~3_combout ;
wire \burst_uncompress_address_base[1]~0_combout ;
wire \burst_uncompress_address_base[1]~q ;
wire \Add2~5_sumout ;
wire \p1_burst_uncompress_address_offset[0]~combout ;
wire \burst_uncompress_address_offset[0]~q ;
wire \Add2~6 ;
wire \Add2~1_sumout ;
wire \p1_burst_uncompress_address_offset[1]~combout ;
wire \burst_uncompress_address_offset[1]~q ;


cyclonev_lcell_comb \last_packet_beat~4 (
	.dataa(!comb),
	.datab(!mem_39_0),
	.datac(!\last_packet_beat~0_combout ),
	.datad(!\last_packet_beat~1_combout ),
	.datae(!\last_packet_beat~2_combout ),
	.dataf(!\last_packet_beat~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~4 .extended_lut = "off";
defparam \last_packet_beat~4 .lut_mask = 64'h3332333233322222;
defparam \last_packet_beat~4 .shared_arith = "off";

cyclonev_lcell_comb \source_addr[1]~0 (
	.dataa(!\burst_uncompress_address_base[1]~q ),
	.datab(!\burst_uncompress_address_offset[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[1]~0 .extended_lut = "off";
defparam \source_addr[1]~0 .lut_mask = 64'h7777777777777777;
defparam \source_addr[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \source_addr[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_94_0),
	.datad(!mem_used_01),
	.datae(!\burst_uncompress_busy~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[1]~1 .extended_lut = "off";
defparam \source_addr[1]~1 .lut_mask = 64'h007F0000007F0000;
defparam \source_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb source_endofpacket(
	.dataa(!mem_95_0),
	.datab(!last_packet_beat),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_endofpacket1),
	.sumout(),
	.cout(),
	.shareout());
defparam source_endofpacket.extended_lut = "off";
defparam source_endofpacket.lut_mask = 64'h4444444444444444;
defparam source_endofpacket.shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!comb),
	.datab(!out_valid),
	.datac(!mem_95_0),
	.datad(!last_packet_beat),
	.datae(!always10),
	.dataf(!p1_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h5155111155555555;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_49_0),
	.datab(!mem_48_0),
	.datac(!mem_47_0),
	.datad(!mem_46_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!\burst_uncompress_byte_counter[2]~q ),
	.datab(!\burst_uncompress_byte_counter[1]~q ),
	.datac(!mem_47_0),
	.datad(!mem_46_0),
	.datae(!last_packet_beat),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000F00F00009999;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \Add0~3 (
	.dataa(!\burst_uncompress_byte_counter[3]~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\burst_uncompress_byte_counter[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~3 .extended_lut = "off";
defparam \Add0~3 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~3 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!mem_48_0),
	.datab(!mem_47_0),
	.datac(!mem_46_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!\burst_uncompress_byte_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \Add1~2 (
	.dataa(!mem_49_0),
	.datab(!mem_48_0),
	.datac(!mem_47_0),
	.datad(!mem_46_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~2 .extended_lut = "off";
defparam \Add1~2 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!last_packet_beat),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~2_combout ),
	.datad(!\Add1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!\burst_uncompress_byte_counter[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAAAAAA6AAAAAAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_50_0),
	.datab(!last_packet_beat),
	.datac(!\burst_uncompress_byte_counter~0_combout ),
	.datad(!\Add1~0_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h1323102013231020;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!\burst_uncompress_byte_counter[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000000080000000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_50_0),
	.datab(!\Add1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h2222222222222222;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!mem_51_0),
	.datac(!last_packet_beat),
	.datad(!\burst_uncompress_byte_counter~0_combout ),
	.datae(!\Add0~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h0305030A0C050C0A;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~7 (
	.dataa(!\burst_uncompress_byte_counter[0]~q ),
	.datab(!\burst_uncompress_busy~q ),
	.datac(!mem_45_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~7 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~7 .lut_mask = 64'h001F0011001F0011;
defparam \burst_uncompress_byte_counter~7 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[0] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[0]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[0] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[0] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(!\burst_uncompress_byte_counter[2]~q ),
	.dataf(!\burst_uncompress_byte_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h8000000000000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~8 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!mem_51_0),
	.datac(!last_packet_beat),
	.datad(!\burst_uncompress_byte_counter~0_combout ),
	.datae(!\Add0~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~8 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~8 .lut_mask = 64'h0000000A0C000C0A;
defparam \burst_uncompress_byte_counter~8 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[1]~q ),
	.datac(!\last_packet_beat~1_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!\last_packet_beat~0_combout ),
	.datab(!mem_46_0),
	.datac(!last_packet_beat),
	.datad(!\burst_uncompress_byte_counter~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h080A080A080A080A;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[1] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_byte_counter[1]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[1] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[1] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h1111111111111111;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_51_0),
	.datac(!mem_50_0),
	.datad(!mem_49_0),
	.datae(!mem_48_0),
	.dataf(!mem_47_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h8000000000000000;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!mem_46_0),
	.datab(!mem_45_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h4444444444444444;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_address_base[1]~0 (
	.dataa(!\burst_uncompress_address_base[1]~q ),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!out_valid1),
	.datae(!p1_ready),
	.dataf(!mem_53_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_address_base[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_address_base[1]~0 .extended_lut = "off";
defparam \burst_uncompress_address_base[1]~0 .lut_mask = 64'h4755474744554444;
defparam \burst_uncompress_address_base[1]~0 .shared_arith = "off";

dffeas \burst_uncompress_address_base[1] (
	.clk(clk),
	.d(\burst_uncompress_address_base[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\burst_uncompress_address_base[1]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_base[1] .is_wysiwyg = "true";
defparam \burst_uncompress_address_base[1] .power_up = "low";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!comb),
	.datab(!\burst_uncompress_busy~q ),
	.datac(!mem_18_0),
	.datad(!mem_59_0),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FB400000FF00;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[0] (
	.dataa(!\Add2~5_sumout ),
	.datab(!mem_52_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[0] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[0] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[0] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[0] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[0]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_address_offset[0]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[0] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[0] .power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!comb),
	.datab(!\burst_uncompress_busy~q ),
	.datac(!mem_19_0),
	.datad(!mem_59_0),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[1]~q ),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FB40000000FF;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[1] (
	.dataa(!mem_53_0),
	.datab(!\Add2~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[1] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[1] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[1] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[1] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[1]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_ready),
	.q(\burst_uncompress_address_offset[1]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[1] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[1] .power_up = "low";

endmodule

module system_altera_merlin_slave_translator (
	WideOr0,
	in_ready_hold,
	read_latency_shift_reg_0,
	m0_write,
	reset,
	in_data_reg_42,
	clk)/* synthesis synthesis_greybox=0 */;
input 	WideOr0;
input 	in_ready_hold;
output 	read_latency_shift_reg_0;
input 	m0_write;
input 	reset;
input 	in_data_reg_42;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!WideOr0),
	.datab(!in_ready_hold),
	.datac(!m0_write),
	.datad(!in_data_reg_42),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module system_altera_merlin_width_adapter (
	h2f_lw_WLAST_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	out_data_49,
	src_data_66,
	saved_grant_1,
	saved_grant_0,
	src_data_78,
	src_data_79,
	src_data_77,
	in_ready,
	nxt_out_eop,
	nxt_out_eop1,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	r_sync_rst,
	use_reg1,
	WideOr1,
	out_endofpacket,
	out_data_59,
	sop_enable,
	address_burst_0,
	out_data_18,
	address_burst_1,
	int_output_sel_0,
	out_data_17,
	out_data_16,
	write_cp_data_69,
	src_payload,
	src_data_69,
	src_data_68,
	Add2,
	src_data_67,
	src_data_65,
	write_cp_data_66,
	src_payload1,
	out_data_50,
	out_data_48,
	ShiftLeft0,
	out_data_47,
	write_cp_data_67,
	out_data_471,
	out_data_51,
	write_cp_data_68,
	src_payload2,
	out_data_511,
	byte_cnt_reg_1,
	out_data_46,
	out_data_461,
	out_data_0,
	address_reg_2,
	src_data_38,
	address_reg_3,
	src_data_39,
	address_reg_4,
	src_payload3,
	out_data_4,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_41,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	in_endofpacket,
	out_data_481,
	out_data_512,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
output 	out_data_49;
input 	src_data_66;
input 	saved_grant_1;
input 	saved_grant_0;
input 	src_data_78;
input 	src_data_79;
input 	src_data_77;
output 	in_ready;
input 	nxt_out_eop;
input 	nxt_out_eop1;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	r_sync_rst;
output 	use_reg1;
input 	WideOr1;
output 	out_endofpacket;
output 	out_data_59;
input 	sop_enable;
input 	address_burst_0;
output 	out_data_18;
input 	address_burst_1;
output 	int_output_sel_0;
output 	out_data_17;
output 	out_data_16;
input 	write_cp_data_69;
input 	src_payload;
input 	src_data_69;
input 	src_data_68;
input 	Add2;
input 	src_data_67;
input 	src_data_65;
input 	write_cp_data_66;
input 	src_payload1;
output 	out_data_50;
output 	out_data_48;
output 	ShiftLeft0;
output 	out_data_47;
input 	write_cp_data_67;
output 	out_data_471;
output 	out_data_51;
input 	write_cp_data_68;
input 	src_payload2;
output 	out_data_511;
output 	byte_cnt_reg_1;
output 	out_data_46;
output 	out_data_461;
output 	out_data_0;
output 	address_reg_2;
input 	src_data_38;
output 	address_reg_3;
input 	src_data_39;
output 	address_reg_4;
input 	src_payload3;
input 	out_data_4;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_41;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
input 	in_endofpacket;
output 	out_data_481;
output 	out_data_512;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add2~0_combout ;
wire \address_reg~0_combout ;
wire \byte_cnt_reg[4]~q ;
wire \Decoder0~0_combout ;
wire \int_byte_cnt_factor[0]~0_combout ;
wire \ShiftLeft0~0_combout ;
wire \Decoder0~1_combout ;
wire \count~0_combout ;
wire \count[0]~1_combout ;
wire \count[0]~q ;
wire \use_reg~0_combout ;
wire \endofpacket_reg~q ;
wire \out_endofpacket~0_combout ;
wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \Decoder0~4_combout ;
wire \LessThan3~0_combout ;
wire \Add1~1_sumout ;
wire \address_reg[0]~q ;
wire \out_data[18]~1_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \address_reg[1]~q ;
wire \int_output_sel[0]~0_combout ;
wire \Add2~1_combout ;
wire \byte_cnt_reg[5]~q ;
wire \out_data[50]~5_combout ;
wire \out_data[50]~6_combout ;
wire \out_data[50]~7_combout ;
wire \Add2~2_combout ;
wire \byte_cnt_reg[3]~q ;
wire \ShiftLeft0~5_combout ;
wire \Add2~3_combout ;
wire \byte_cnt_reg[2]~q ;
wire \out_data[47]~11_combout ;
wire \ShiftLeft0~2_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \Add2~4_combout ;
wire \byte_cnt_reg[6]~q ;
wire \out_data[51]~14_combout ;
wire \byte_cnt_reg~0_combout ;
wire \Decoder0~5_combout ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \Decoder0~6_combout ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add1~14 ;
wire \Add1~17_sumout ;


cyclonev_lcell_comb \out_data[49]~36 (
	.dataa(!src_data_65),
	.datab(!src_data_77),
	.datac(!\byte_cnt_reg[4]~q ),
	.datad(!src_data_78),
	.datae(!use_reg1),
	.dataf(!\ShiftLeft0~0_combout ),
	.datag(!src_data_79),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[49]~36 .extended_lut = "on";
defparam \out_data[49]~36 .lut_mask = 64'h04000F0FF4F00F0F;
defparam \out_data[49]~36 .shared_arith = "off";

cyclonev_lcell_comb \in_ready~0 (
	.dataa(!saved_grant_1),
	.datab(!\count[0]~q ),
	.datac(!src_data_78),
	.datad(!src_data_79),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_ready~0 .extended_lut = "off";
defparam \in_ready~0 .lut_mask = 64'h0888088808880888;
defparam \in_ready~0 .shared_arith = "off";

dffeas use_reg(
	.clk(clk_clk),
	.d(\use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(use_reg1),
	.prn(vcc));
defparam use_reg.is_wysiwyg = "true";
defparam use_reg.power_up = "low";

cyclonev_lcell_comb \out_endofpacket~1 (
	.dataa(!saved_grant_1),
	.datab(!\count[0]~q ),
	.datac(!use_reg1),
	.datad(!\endofpacket_reg~q ),
	.datae(!\out_endofpacket~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_endofpacket),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~1 .extended_lut = "off";
defparam \out_endofpacket~1 .lut_mask = 64'h5457FCFF5457FCFF;
defparam \out_endofpacket~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[59]~0 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_59),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[59]~0 .extended_lut = "off";
defparam \out_data[59]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \out_data[59]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[18]~2 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(gnd),
	.datad(!use_reg1),
	.datae(!\address_reg[0]~q ),
	.dataf(!\out_data[18]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[18]~2 .extended_lut = "off";
defparam \out_data[18]~2 .lut_mask = 64'h000000FF880088FF;
defparam \out_data[18]~2 .shared_arith = "off";

cyclonev_lcell_comb \int_output_sel[0]~1 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(gnd),
	.datad(!use_reg1),
	.datae(!\address_reg[1]~q ),
	.dataf(!\int_output_sel[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(int_output_sel_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[0]~1 .extended_lut = "off";
defparam \int_output_sel[0]~1 .lut_mask = 64'h000000FF880088FF;
defparam \int_output_sel[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[17]~3 (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!h2f_lw_WSTRB_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[17]~3 .extended_lut = "off";
defparam \out_data[17]~3 .lut_mask = 64'h0F5F0F3F0F5F0F3F;
defparam \out_data[17]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[16]~4 (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!h2f_lw_WSTRB_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[16]~4 .extended_lut = "off";
defparam \out_data[16]~4 .lut_mask = 64'h0F5F0F3F0F5F0F3F;
defparam \out_data[16]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[50]~8 (
	.dataa(!src_data_78),
	.datab(!use_reg1),
	.datac(!\byte_cnt_reg[5]~q ),
	.datad(!\out_data[50]~5_combout ),
	.datae(!\out_data[50]~6_combout ),
	.dataf(!\out_data[50]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[50]~8 .extended_lut = "off";
defparam \out_data[50]~8 .lut_mask = 64'h03FF8BFF8BFF8BFF;
defparam \out_data[50]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_data[48]~9 (
	.dataa(!use_reg1),
	.datab(!\byte_cnt_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[48]~9 .extended_lut = "off";
defparam \out_data[48]~9 .lut_mask = 64'h1111111111111111;
defparam \out_data[48]~9 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!src_data_68),
	.datab(!src_data_67),
	.datac(!src_data_66),
	.datad(!src_data_65),
	.datae(!\int_byte_cnt_factor[0]~0_combout ),
	.dataf(!src_data_78),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h3333555500FF0F0F;
defparam \ShiftLeft0~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[47]~10 (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!use_reg1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[47]~10 .extended_lut = "off";
defparam \out_data[47]~10 .lut_mask = 64'hFAC80000FAC80000;
defparam \out_data[47]~10 .shared_arith = "off";

cyclonev_lcell_comb \out_data[47]~12 (
	.dataa(!src_data_78),
	.datab(!out_data_47),
	.datac(!\out_data[47]~11_combout ),
	.datad(!\ShiftLeft0~2_combout ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\ShiftLeft0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_471),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[47]~12 .extended_lut = "off";
defparam \out_data[47]~12 .lut_mask = 64'h0F2F2F2F3F3F3F3F;
defparam \out_data[47]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_data[51]~13 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!use_reg1),
	.datad(!\ShiftLeft0~2_combout ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\ShiftLeft0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[51]~13 .extended_lut = "off";
defparam \out_data[51]~13 .lut_mask = 64'h0020202030303030;
defparam \out_data[51]~13 .shared_arith = "off";

cyclonev_lcell_comb \out_data[51]~15 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!use_reg1),
	.datad(!\byte_cnt_reg[6]~q ),
	.datae(!\out_data[51]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_511),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[51]~15 .extended_lut = "off";
defparam \out_data[51]~15 .lut_mask = 64'h404F000F404F000F;
defparam \out_data[51]~15 .shared_arith = "off";

dffeas \byte_cnt_reg[1] (
	.clk(clk_clk),
	.d(\byte_cnt_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(byte_cnt_reg_1),
	.prn(vcc));
defparam \byte_cnt_reg[1] .is_wysiwyg = "true";
defparam \byte_cnt_reg[1] .power_up = "low";

cyclonev_lcell_comb \out_data[46]~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\Decoder0~0_combout ),
	.datad(!src_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[46]~16 .extended_lut = "off";
defparam \out_data[46]~16 .lut_mask = 64'h000F000F000F000F;
defparam \out_data[46]~16 .shared_arith = "off";

cyclonev_lcell_comb \out_data[46]~17 (
	.dataa(gnd),
	.datab(!use_reg1),
	.datac(!\Decoder0~0_combout ),
	.datad(!byte_cnt_reg_1),
	.datae(!src_data_65),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_461),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[46]~17 .extended_lut = "off";
defparam \out_data[46]~17 .lut_mask = 64'h00330C3F00330C3F;
defparam \out_data[46]~17 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~18 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!h2f_lw_WDATA_16),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~18 .extended_lut = "off";
defparam \out_data[0]~18 .lut_mask = 64'h5353535353535353;
defparam \out_data[0]~18 .shared_arith = "off";

dffeas \address_reg[2] (
	.clk(clk_clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_2),
	.prn(vcc));
defparam \address_reg[2] .is_wysiwyg = "true";
defparam \address_reg[2] .power_up = "low";

dffeas \address_reg[3] (
	.clk(clk_clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_3),
	.prn(vcc));
defparam \address_reg[3] .is_wysiwyg = "true";
defparam \address_reg[3] .power_up = "low";

dffeas \address_reg[4] (
	.clk(clk_clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_4),
	.prn(vcc));
defparam \address_reg[4] .is_wysiwyg = "true";
defparam \address_reg[4] .power_up = "low";

cyclonev_lcell_comb \out_data[1]~19 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!h2f_lw_WDATA_17),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~19 .extended_lut = "off";
defparam \out_data[1]~19 .lut_mask = 64'h5353535353535353;
defparam \out_data[1]~19 .shared_arith = "off";

cyclonev_lcell_comb \out_data[2]~20 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!h2f_lw_WDATA_18),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~20 .extended_lut = "off";
defparam \out_data[2]~20 .lut_mask = 64'h5353535353535353;
defparam \out_data[2]~20 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~21 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!h2f_lw_WDATA_19),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~21 .extended_lut = "off";
defparam \out_data[3]~21 .lut_mask = 64'h5353535353535353;
defparam \out_data[3]~21 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~22 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!h2f_lw_WDATA_20),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~22 .extended_lut = "off";
defparam \out_data[4]~22 .lut_mask = 64'h5353535353535353;
defparam \out_data[4]~22 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~23 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!h2f_lw_WDATA_21),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~23 .extended_lut = "off";
defparam \out_data[5]~23 .lut_mask = 64'h5353535353535353;
defparam \out_data[5]~23 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~24 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!h2f_lw_WDATA_22),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~24 .extended_lut = "off";
defparam \out_data[6]~24 .lut_mask = 64'h5353535353535353;
defparam \out_data[6]~24 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~25 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!h2f_lw_WDATA_23),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~25 .extended_lut = "off";
defparam \out_data[7]~25 .lut_mask = 64'h5353535353535353;
defparam \out_data[7]~25 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~26 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!h2f_lw_WDATA_24),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~26 .extended_lut = "off";
defparam \out_data[8]~26 .lut_mask = 64'h5353535353535353;
defparam \out_data[8]~26 .shared_arith = "off";

cyclonev_lcell_comb \out_data[9]~27 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!h2f_lw_WDATA_25),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[9]~27 .extended_lut = "off";
defparam \out_data[9]~27 .lut_mask = 64'h5353535353535353;
defparam \out_data[9]~27 .shared_arith = "off";

cyclonev_lcell_comb \out_data[10]~28 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!h2f_lw_WDATA_26),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[10]~28 .extended_lut = "off";
defparam \out_data[10]~28 .lut_mask = 64'h5353535353535353;
defparam \out_data[10]~28 .shared_arith = "off";

cyclonev_lcell_comb \out_data[11]~29 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!h2f_lw_WDATA_27),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[11]~29 .extended_lut = "off";
defparam \out_data[11]~29 .lut_mask = 64'h5353535353535353;
defparam \out_data[11]~29 .shared_arith = "off";

cyclonev_lcell_comb \out_data[12]~30 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!h2f_lw_WDATA_28),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[12]~30 .extended_lut = "off";
defparam \out_data[12]~30 .lut_mask = 64'h5353535353535353;
defparam \out_data[12]~30 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~31 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!h2f_lw_WDATA_29),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~31 .extended_lut = "off";
defparam \out_data[13]~31 .lut_mask = 64'h5353535353535353;
defparam \out_data[13]~31 .shared_arith = "off";

cyclonev_lcell_comb \out_data[14]~32 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!h2f_lw_WDATA_30),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[14]~32 .extended_lut = "off";
defparam \out_data[14]~32 .lut_mask = 64'h5353535353535353;
defparam \out_data[14]~32 .shared_arith = "off";

cyclonev_lcell_comb \out_data[15]~33 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!h2f_lw_WDATA_31),
	.datac(!int_output_sel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[15]~33 .extended_lut = "off";
defparam \out_data[15]~33 .lut_mask = 64'h5353535353535353;
defparam \out_data[15]~33 .shared_arith = "off";

cyclonev_lcell_comb \out_data[48]~34 (
	.dataa(!out_data_48),
	.datab(!ShiftLeft0),
	.datac(!out_data_47),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_481),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[48]~34 .extended_lut = "off";
defparam \out_data[48]~34 .lut_mask = 64'h5757575757575757;
defparam \out_data[48]~34 .shared_arith = "off";

cyclonev_lcell_comb \out_data[51]~35 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!use_reg1),
	.datad(!\ShiftLeft0~5_combout ),
	.datae(!\byte_cnt_reg[6]~q ),
	.dataf(!\out_data[51]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_512),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[51]~35 .extended_lut = "off";
defparam \out_data[51]~35 .lut_mask = 64'h40704F7F00300F3F;
defparam \out_data[51]~35 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!out_data_461),
	.datab(!out_data_481),
	.datac(!out_data_471),
	.datad(!out_data_49),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h807F807F807F807F;
defparam \Add2~0 .shared_arith = "off";

cyclonev_lcell_comb \address_reg~0 (
	.dataa(!nxt_out_eop),
	.datab(!nxt_out_eop1),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(!use_reg1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_reg~0 .extended_lut = "off";
defparam \address_reg~0 .lut_mask = 64'hFFFFFF07FFFFFF07;
defparam \address_reg~0 .shared_arith = "off";

dffeas \byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\Add2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[4]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \byte_cnt_reg[4] .power_up = "low";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!h2f_lw_AWSIZE_1),
	.datad(!h2f_lw_AWSIZE_2),
	.datae(!saved_grant_1),
	.dataf(!saved_grant_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'hFFFF8888F0008000;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \int_byte_cnt_factor[0]~0 (
	.dataa(!src_data_77),
	.datab(!\Decoder0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_byte_cnt_factor[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_byte_cnt_factor[0]~0 .extended_lut = "off";
defparam \int_byte_cnt_factor[0]~0 .lut_mask = 64'h8888888888888888;
defparam \int_byte_cnt_factor[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!src_data_69),
	.datab(!src_data_68),
	.datac(!src_data_67),
	.datad(!src_data_66),
	.datae(!\int_byte_cnt_factor[0]~0_combout ),
	.dataf(!src_data_78),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h3333AAAA00FF0F0F;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!src_data_77),
	.datab(!\Decoder0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h1111111111111111;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \count~0 (
	.dataa(!saved_grant_1),
	.datab(!src_data_78),
	.datac(!src_data_79),
	.datad(gnd),
	.datae(!WideOr1),
	.dataf(!use_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~0 .extended_lut = "off";
defparam \count~0 .lut_mask = 64'h00002A2A00000000;
defparam \count~0 .shared_arith = "off";

cyclonev_lcell_comb \count[0]~1 (
	.dataa(!\count[0]~q ),
	.datab(!nxt_in_ready2),
	.datac(!nxt_in_ready1),
	.datad(!use_reg1),
	.datae(!\Decoder0~1_combout ),
	.dataf(!\count~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[0]~1 .extended_lut = "off";
defparam \count[0]~1 .lut_mask = 64'h55A655A6F7A604A6;
defparam \count[0]~1 .shared_arith = "off";

dffeas \count[0] (
	.clk(clk_clk),
	.d(\count[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclonev_lcell_comb \use_reg~0 (
	.dataa(!\count[0]~q ),
	.datab(!nxt_in_ready2),
	.datac(!nxt_in_ready1),
	.datad(!use_reg1),
	.datae(!\count~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\use_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \use_reg~0 .extended_lut = "off";
defparam \use_reg~0 .lut_mask = 64'h00AEF3FF00AEF3FF;
defparam \use_reg~0 .shared_arith = "off";

dffeas endofpacket_reg(
	.clk(clk_clk),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!use_reg1),
	.q(\endofpacket_reg~q ),
	.prn(vcc));
defparam endofpacket_reg.is_wysiwyg = "true";
defparam endofpacket_reg.power_up = "low";

cyclonev_lcell_comb \out_endofpacket~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_0),
	.datac(!src_data_78),
	.datad(!src_data_79),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_endofpacket~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~0 .extended_lut = "off";
defparam \out_endofpacket~0 .lut_mask = 64'h1000100010001000;
defparam \out_endofpacket~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!src_data_77),
	.datab(!\Decoder0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h2222222222222222;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h6E6E6E6E6E6E6E6E;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\Decoder0~2_combout ),
	.datab(!\Decoder0~3_combout ),
	.datac(!\Decoder0~4_combout ),
	.datad(!out_data_18),
	.datae(gnd),
	.dataf(!\LessThan3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000F7FF000000FF;
defparam \Add1~1 .shared_arith = "off";

dffeas \address_reg[0] (
	.clk(clk_clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[0]~q ),
	.prn(vcc));
defparam \address_reg[0] .is_wysiwyg = "true";
defparam \address_reg[0] .power_up = "low";

cyclonev_lcell_comb \out_data[18]~1 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!h2f_lw_AWADDR_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!address_burst_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[18]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[18]~1 .extended_lut = "off";
defparam \out_data[18]~1 .lut_mask = 64'h05370505053705FF;
defparam \out_data[18]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!\Decoder0~2_combout ),
	.datab(!\Decoder0~3_combout ),
	.datac(!\Decoder0~1_combout ),
	.datad(!int_output_sel_0),
	.datae(gnd),
	.dataf(!\LessThan3~0_combout ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h00008000000000FF;
defparam \Add1~5 .shared_arith = "off";

dffeas \address_reg[1] (
	.clk(clk_clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[1]~q ),
	.prn(vcc));
defparam \address_reg[1] .is_wysiwyg = "true";
defparam \address_reg[1] .power_up = "low";

cyclonev_lcell_comb \int_output_sel[0]~0 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!h2f_lw_AWADDR_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!address_burst_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_output_sel[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[0]~0 .extended_lut = "off";
defparam \int_output_sel[0]~0 .lut_mask = 64'h05370505053705FF;
defparam \int_output_sel[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!out_data_461),
	.datab(!out_data_481),
	.datac(!out_data_471),
	.datad(!out_data_49),
	.datae(!out_data_50),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h80007FFF80007FFF;
defparam \Add2~1 .shared_arith = "off";

dffeas \byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\Add2~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[5]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \byte_cnt_reg[5] .power_up = "low";

cyclonev_lcell_comb \out_data[50]~5 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(!use_reg1),
	.datae(!src_data_68),
	.dataf(!src_data_67),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[50]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[50]~5 .extended_lut = "off";
defparam \out_data[50]~5 .lut_mask = 64'h0000400004004400;
defparam \out_data[50]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[50]~6 (
	.dataa(!saved_grant_0),
	.datab(!src_data_78),
	.datac(!src_data_79),
	.datad(!src_data_77),
	.datae(!write_cp_data_69),
	.dataf(!src_payload),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[50]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[50]~6 .extended_lut = "off";
defparam \out_data[50]~6 .lut_mask = 64'h00004050C0F0C0F0;
defparam \out_data[50]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[50]~7 (
	.dataa(!saved_grant_0),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(!src_data_65),
	.datae(!write_cp_data_66),
	.dataf(!src_payload1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[50]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[50]~7 .extended_lut = "off";
defparam \out_data[50]~7 .lut_mask = 64'h0003101330333033;
defparam \out_data[50]~7 .shared_arith = "off";

cyclonev_lcell_comb \Add2~2 (
	.dataa(!out_data_461),
	.datab(!out_data_48),
	.datac(!ShiftLeft0),
	.datad(!out_data_47),
	.datae(!out_data_471),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~2 .extended_lut = "off";
defparam \Add2~2 .lut_mask = 64'h9995333F9995333F;
defparam \Add2~2 .shared_arith = "off";

dffeas \byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\Add2~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[3]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \byte_cnt_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(!src_data_65),
	.datae(!src_data_66),
	.dataf(!src_data_67),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "off";
defparam \ShiftLeft0~5 .lut_mask = 64'h00508ADA2070AAFA;
defparam \ShiftLeft0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add2~3 (
	.dataa(!out_data_461),
	.datab(!out_data_47),
	.datac(!\out_data[47]~11_combout ),
	.datad(!\ShiftLeft0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~3 .extended_lut = "off";
defparam \Add2~3 .lut_mask = 64'hA595A595A595A595;
defparam \Add2~3 .shared_arith = "off";

dffeas \byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\Add2~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[2]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \byte_cnt_reg[2] .power_up = "low";

cyclonev_lcell_comb \out_data[47]~11 (
	.dataa(!use_reg1),
	.datab(!\byte_cnt_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[47]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[47]~11 .extended_lut = "off";
defparam \out_data[47]~11 .lut_mask = 64'h1111111111111111;
defparam \out_data[47]~11 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!src_data_77),
	.datad(!\Decoder0~0_combout ),
	.datae(!write_cp_data_67),
	.dataf(!Add2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h0000300050007000;
defparam \ShiftLeft0~2 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!saved_grant_0),
	.datab(!src_data_77),
	.datac(!\Decoder0~0_combout ),
	.datad(!write_cp_data_66),
	.datae(!src_payload1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h00153F3F00153F3F;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!src_data_78),
	.datab(gnd),
	.datac(!src_data_77),
	.datad(!src_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h0050005000500050;
defparam \ShiftLeft0~4 .shared_arith = "off";

cyclonev_lcell_comb \Add2~4 (
	.dataa(!out_data_461),
	.datab(!out_data_481),
	.datac(!out_data_471),
	.datad(!out_data_49),
	.datae(!out_data_50),
	.dataf(!out_data_512),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~4 .extended_lut = "off";
defparam \Add2~4 .lut_mask = 64'h800000007FFFFFFF;
defparam \Add2~4 .shared_arith = "off";

dffeas \byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\Add2~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[6]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \byte_cnt_reg[6] .power_up = "low";

cyclonev_lcell_comb \out_data[51]~14 (
	.dataa(!saved_grant_0),
	.datab(!src_data_77),
	.datac(!write_cp_data_68),
	.datad(!src_payload2),
	.datae(!write_cp_data_69),
	.dataf(!src_payload),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[51]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[51]~14 .extended_lut = "off";
defparam \out_data[51]~14 .lut_mask = 64'hFECCBA8832003200;
defparam \out_data[51]~14 .shared_arith = "off";

cyclonev_lcell_comb \byte_cnt_reg~0 (
	.dataa(!nxt_in_ready2),
	.datab(!nxt_in_ready1),
	.datac(!use_reg1),
	.datad(!byte_cnt_reg_1),
	.datae(!out_data_46),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_cnt_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_cnt_reg~0 .extended_lut = "off";
defparam \byte_cnt_reg~0 .lut_mask = 64'hFDF20D02FDF20D02;
defparam \byte_cnt_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!use_reg1),
	.datab(!out_data_59),
	.datac(!\Decoder0~5_combout ),
	.datad(!address_reg_2),
	.datae(gnd),
	.dataf(!src_data_38),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FB510000085D;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~6 (
	.dataa(!src_data_78),
	.datab(!src_data_79),
	.datac(!src_data_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~6 .extended_lut = "off";
defparam \Decoder0~6 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~6 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!use_reg1),
	.datab(!out_data_59),
	.datac(!\Decoder0~6_combout ),
	.datad(!address_reg_3),
	.datae(gnd),
	.dataf(!src_data_39),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FB510000085D;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!saved_grant_0),
	.datab(!use_reg1),
	.datac(!out_data_4),
	.datad(!src_payload3),
	.datae(gnd),
	.dataf(!address_reg_4),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFCC000004CC;
defparam \Add1~17 .shared_arith = "off";

endmodule

module system_altera_merlin_width_adapter_1 (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	always10,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_94_0,
	mem_used_01,
	out_valid,
	mem_95_0,
	mem_39_0,
	last_packet_beat,
	source_addr_1,
	source_addr_11,
	mem_19_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_59_0,
	mem_41_0,
	mem_0_0,
	out_data_0,
	mem_1_0,
	out_data_1,
	mem_2_0,
	out_data_2,
	mem_3_0,
	out_data_3,
	mem_4_0,
	out_data_4,
	mem_5_0,
	out_data_5,
	mem_6_0,
	out_data_6,
	mem_7_0,
	out_data_7,
	mem_8_0,
	out_data_8,
	mem_9_0,
	out_data_9,
	mem_10_0,
	out_data_10,
	mem_11_0,
	out_data_11,
	mem_12_0,
	out_data_12,
	mem_13_0,
	out_data_13,
	mem_14_0,
	out_data_14,
	mem_15_0,
	out_data_15,
	ShiftLeft2,
	ShiftLeft21,
	ShiftLeft22,
	ShiftLeft23,
	ShiftLeft24,
	ShiftLeft25,
	ShiftLeft26,
	ShiftLeft27,
	ShiftLeft28,
	ShiftLeft29,
	ShiftLeft210,
	ShiftLeft211,
	ShiftLeft212,
	ShiftLeft213,
	ShiftLeft214,
	ShiftLeft215,
	r_sync_rst,
	p1_ready,
	out_valid1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
output 	always10;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_94_0;
input 	mem_used_01;
output 	out_valid;
input 	mem_95_0;
input 	mem_39_0;
input 	last_packet_beat;
input 	source_addr_1;
input 	source_addr_11;
input 	mem_19_0;
input 	mem_91_0;
input 	mem_92_0;
input 	mem_93_0;
input 	mem_59_0;
input 	mem_41_0;
input 	mem_0_0;
output 	out_data_0;
input 	mem_1_0;
output 	out_data_1;
input 	mem_2_0;
output 	out_data_2;
input 	mem_3_0;
output 	out_data_3;
input 	mem_4_0;
output 	out_data_4;
input 	mem_5_0;
output 	out_data_5;
input 	mem_6_0;
output 	out_data_6;
input 	mem_7_0;
output 	out_data_7;
input 	mem_8_0;
output 	out_data_8;
input 	mem_9_0;
output 	out_data_9;
input 	mem_10_0;
output 	out_data_10;
input 	mem_11_0;
output 	out_data_11;
input 	mem_12_0;
output 	out_data_12;
input 	mem_13_0;
output 	out_data_13;
input 	mem_14_0;
output 	out_data_14;
input 	mem_15_0;
output 	out_data_15;
output 	ShiftLeft2;
output 	ShiftLeft21;
output 	ShiftLeft22;
output 	ShiftLeft23;
output 	ShiftLeft24;
output 	ShiftLeft25;
output 	ShiftLeft26;
output 	ShiftLeft27;
output 	ShiftLeft28;
output 	ShiftLeft29;
output 	ShiftLeft210;
output 	ShiftLeft211;
output 	ShiftLeft212;
output 	ShiftLeft213;
output 	ShiftLeft214;
output 	ShiftLeft215;
input 	r_sync_rst;
output 	p1_ready;
output 	out_valid1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ShiftLeft2~0_combout ;
wire \data_reg~0_combout ;
wire \always10~0_combout ;
wire \always9~0_combout ;
wire \data_reg[0]~q ;
wire \LessThan13~0_combout ;
wire \ShiftLeft2~1_combout ;
wire \data_reg~1_combout ;
wire \data_reg[1]~q ;
wire \ShiftLeft2~2_combout ;
wire \data_reg~2_combout ;
wire \data_reg[2]~q ;
wire \ShiftLeft2~3_combout ;
wire \data_reg~3_combout ;
wire \data_reg[3]~q ;
wire \ShiftLeft2~4_combout ;
wire \data_reg~4_combout ;
wire \data_reg[4]~q ;
wire \ShiftLeft2~5_combout ;
wire \data_reg~5_combout ;
wire \data_reg[5]~q ;
wire \ShiftLeft2~6_combout ;
wire \data_reg~6_combout ;
wire \data_reg[6]~q ;
wire \ShiftLeft2~7_combout ;
wire \data_reg~7_combout ;
wire \data_reg[7]~q ;
wire \ShiftLeft2~8_combout ;
wire \data_reg~8_combout ;
wire \data_reg[8]~q ;
wire \ShiftLeft2~9_combout ;
wire \data_reg~9_combout ;
wire \data_reg[9]~q ;
wire \ShiftLeft2~10_combout ;
wire \data_reg~10_combout ;
wire \data_reg[10]~q ;
wire \ShiftLeft2~11_combout ;
wire \data_reg~11_combout ;
wire \data_reg[11]~q ;
wire \ShiftLeft2~12_combout ;
wire \data_reg~12_combout ;
wire \data_reg[12]~q ;
wire \ShiftLeft2~13_combout ;
wire \data_reg~13_combout ;
wire \data_reg[13]~q ;
wire \ShiftLeft2~14_combout ;
wire \data_reg~14_combout ;
wire \data_reg[14]~q ;
wire \ShiftLeft2~15_combout ;
wire \data_reg~15_combout ;
wire \data_reg[15]~q ;


cyclonev_lcell_comb \always10~1 (
	.dataa(!mem_59_0),
	.datab(!mem_93_0),
	.datac(!mem_19_0),
	.datad(!mem_92_0),
	.datae(!source_addr_11),
	.dataf(!mem_91_0),
	.datag(!source_addr_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(always10),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "on";
defparam \always10~1 .lut_mask = 64'hCF0FCF0F4F0F4F0F;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \out_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_94_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_valid~0 .extended_lut = "off";
defparam \out_valid~0 .lut_mask = 64'h8880888088808880;
defparam \out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~0 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[0]~q ),
	.datae(!\LessThan13~0_combout ),
	.dataf(!\ShiftLeft2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~0 .extended_lut = "off";
defparam \out_data[0]~0 .lut_mask = 64'h00FF0000B8FFB8B8;
defparam \out_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~1 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[1]~q ),
	.dataf(!\ShiftLeft2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~1 .extended_lut = "off";
defparam \out_data[1]~1 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[2]~2 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[2]~q ),
	.dataf(!\ShiftLeft2~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~2 .extended_lut = "off";
defparam \out_data[2]~2 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~3 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[3]~q ),
	.dataf(!\ShiftLeft2~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~3 .extended_lut = "off";
defparam \out_data[3]~3 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~4 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[4]~q ),
	.dataf(!\ShiftLeft2~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~4 .extended_lut = "off";
defparam \out_data[4]~4 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~5 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[5]~q ),
	.dataf(!\ShiftLeft2~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~5 .extended_lut = "off";
defparam \out_data[5]~5 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~6 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[6]~q ),
	.dataf(!\ShiftLeft2~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~6 .extended_lut = "off";
defparam \out_data[6]~6 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~7 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[7]~q ),
	.dataf(!\ShiftLeft2~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~7 .extended_lut = "off";
defparam \out_data[7]~7 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~8 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[8]~q ),
	.dataf(!\ShiftLeft2~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~8 .extended_lut = "off";
defparam \out_data[8]~8 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_data[9]~9 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[9]~q ),
	.dataf(!\ShiftLeft2~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[9]~9 .extended_lut = "off";
defparam \out_data[9]~9 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[9]~9 .shared_arith = "off";

cyclonev_lcell_comb \out_data[10]~10 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[10]~q ),
	.dataf(!\ShiftLeft2~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[10]~10 .extended_lut = "off";
defparam \out_data[10]~10 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[10]~10 .shared_arith = "off";

cyclonev_lcell_comb \out_data[11]~11 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[11]~q ),
	.dataf(!\ShiftLeft2~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[11]~11 .extended_lut = "off";
defparam \out_data[11]~11 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[11]~11 .shared_arith = "off";

cyclonev_lcell_comb \out_data[12]~12 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[12]~q ),
	.dataf(!\ShiftLeft2~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[12]~12 .extended_lut = "off";
defparam \out_data[12]~12 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~13 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[13]~q ),
	.dataf(!\ShiftLeft2~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~13 .extended_lut = "off";
defparam \out_data[13]~13 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[13]~13 .shared_arith = "off";

cyclonev_lcell_comb \out_data[14]~14 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[14]~q ),
	.dataf(!\ShiftLeft2~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[14]~14 .extended_lut = "off";
defparam \out_data[14]~14 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[14]~14 .shared_arith = "off";

cyclonev_lcell_comb \out_data[15]~15 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\LessThan13~0_combout ),
	.datae(!\data_reg[15]~q ),
	.dataf(!\ShiftLeft2~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[15]~15 .extended_lut = "off";
defparam \out_data[15]~15 .lut_mask = 64'h0000FF00B8B8FFB8;
defparam \out_data[15]~15 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~16 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft2),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~16 .extended_lut = "off";
defparam \ShiftLeft2~16 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~16 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~17 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft21),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~17 .extended_lut = "off";
defparam \ShiftLeft2~17 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~17 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~18 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft22),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~18 .extended_lut = "off";
defparam \ShiftLeft2~18 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~18 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~19 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft23),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~19 .extended_lut = "off";
defparam \ShiftLeft2~19 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~19 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~20 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft24),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~20 .extended_lut = "off";
defparam \ShiftLeft2~20 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~20 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~21 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft25),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~21 .extended_lut = "off";
defparam \ShiftLeft2~21 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~21 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~22 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft26),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~22 .extended_lut = "off";
defparam \ShiftLeft2~22 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~22 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~23 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft27),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~23 .extended_lut = "off";
defparam \ShiftLeft2~23 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~23 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~24 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft28),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~24 .extended_lut = "off";
defparam \ShiftLeft2~24 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~24 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~25 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft29),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~25 .extended_lut = "off";
defparam \ShiftLeft2~25 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~25 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~26 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft210),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~26 .extended_lut = "off";
defparam \ShiftLeft2~26 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~26 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~27 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft211),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~27 .extended_lut = "off";
defparam \ShiftLeft2~27 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~27 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~28 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~12_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft212),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~28 .extended_lut = "off";
defparam \ShiftLeft2~28 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~28 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~29 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~13_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft213),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~29 .extended_lut = "off";
defparam \ShiftLeft2~29 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~29 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~30 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft214),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~30 .extended_lut = "off";
defparam \ShiftLeft2~30 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~30 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~31 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\ShiftLeft2~15_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft215),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~31 .extended_lut = "off";
defparam \ShiftLeft2~31 .lut_mask = 64'h0047004700470047;
defparam \ShiftLeft2~31 .shared_arith = "off";

cyclonev_lcell_comb \p1_ready~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_39_0),
	.datad(!mem_41_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(p1_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_ready~0 .extended_lut = "off";
defparam \p1_ready~0 .lut_mask = 64'h3353335333533353;
defparam \p1_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \out_valid~1 (
	.dataa(!out_valid),
	.datab(!mem_95_0),
	.datac(!last_packet_beat),
	.datad(!always10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_valid~1 .extended_lut = "off";
defparam \out_valid~1 .lut_mask = 64'h20AA20AA20AA20AA;
defparam \out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~0 (
	.dataa(!q_a_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_0_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~0 .extended_lut = "off";
defparam \ShiftLeft2~0 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~0 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~0 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[0]~q ),
	.datae(!\ShiftLeft2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~0 .extended_lut = "off";
defparam \data_reg~0 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!mem_95_0),
	.datab(!last_packet_beat),
	.datac(!always10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'h4F4F4F4F4F4F4F4F;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \always9~0 (
	.dataa(!out_valid),
	.datab(!mem_95_0),
	.datac(!last_packet_beat),
	.datad(!always10),
	.datae(!p1_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'h8A00AAAA8A00AAAA;
defparam \always9~0 .shared_arith = "off";

dffeas \data_reg[0] (
	.clk(clk_clk),
	.d(\data_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[0]~q ),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

cyclonev_lcell_comb \LessThan13~0 (
	.dataa(!mem_92_0),
	.datab(!mem_91_0),
	.datac(!mem_93_0),
	.datad(!mem_59_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan13~0 .extended_lut = "off";
defparam \LessThan13~0 .lut_mask = 64'h80A080A080A080A0;
defparam \LessThan13~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft2~1 (
	.dataa(!q_a_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_1_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~1 .extended_lut = "off";
defparam \ShiftLeft2~1 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~1 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~1 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[1]~q ),
	.datae(!\ShiftLeft2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~1 .extended_lut = "off";
defparam \data_reg~1 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~1 .shared_arith = "off";

dffeas \data_reg[1] (
	.clk(clk_clk),
	.d(\data_reg~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[1]~q ),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~2 (
	.dataa(!q_a_2),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_2_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~2 .extended_lut = "off";
defparam \ShiftLeft2~2 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~2 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~2 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[2]~q ),
	.datae(!\ShiftLeft2~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~2 .extended_lut = "off";
defparam \data_reg~2 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~2 .shared_arith = "off";

dffeas \data_reg[2] (
	.clk(clk_clk),
	.d(\data_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[2]~q ),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~3 (
	.dataa(!q_a_3),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_3_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~3 .extended_lut = "off";
defparam \ShiftLeft2~3 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~3 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~3 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[3]~q ),
	.datae(!\ShiftLeft2~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~3 .extended_lut = "off";
defparam \data_reg~3 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~3 .shared_arith = "off";

dffeas \data_reg[3] (
	.clk(clk_clk),
	.d(\data_reg~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[3]~q ),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~4 (
	.dataa(!q_a_4),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_4_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~4 .extended_lut = "off";
defparam \ShiftLeft2~4 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~4 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~4 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[4]~q ),
	.datae(!\ShiftLeft2~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~4 .extended_lut = "off";
defparam \data_reg~4 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~4 .shared_arith = "off";

dffeas \data_reg[4] (
	.clk(clk_clk),
	.d(\data_reg~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[4]~q ),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~5 (
	.dataa(!q_a_5),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_5_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~5 .extended_lut = "off";
defparam \ShiftLeft2~5 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~5 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~5 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[5]~q ),
	.datae(!\ShiftLeft2~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~5 .extended_lut = "off";
defparam \data_reg~5 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~5 .shared_arith = "off";

dffeas \data_reg[5] (
	.clk(clk_clk),
	.d(\data_reg~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[5]~q ),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~6 (
	.dataa(!q_a_6),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_6_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~6 .extended_lut = "off";
defparam \ShiftLeft2~6 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~6 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~6 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[6]~q ),
	.datae(!\ShiftLeft2~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~6 .extended_lut = "off";
defparam \data_reg~6 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~6 .shared_arith = "off";

dffeas \data_reg[6] (
	.clk(clk_clk),
	.d(\data_reg~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[6]~q ),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~7 (
	.dataa(!q_a_7),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_7_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~7 .extended_lut = "off";
defparam \ShiftLeft2~7 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~7 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~7 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[7]~q ),
	.datae(!\ShiftLeft2~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~7 .extended_lut = "off";
defparam \data_reg~7 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~7 .shared_arith = "off";

dffeas \data_reg[7] (
	.clk(clk_clk),
	.d(\data_reg~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[7]~q ),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~8 (
	.dataa(!q_a_8),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_8_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~8 .extended_lut = "off";
defparam \ShiftLeft2~8 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~8 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~8 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[8]~q ),
	.datae(!\ShiftLeft2~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~8 .extended_lut = "off";
defparam \data_reg~8 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~8 .shared_arith = "off";

dffeas \data_reg[8] (
	.clk(clk_clk),
	.d(\data_reg~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[8]~q ),
	.prn(vcc));
defparam \data_reg[8] .is_wysiwyg = "true";
defparam \data_reg[8] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~9 (
	.dataa(!q_a_9),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_9_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~9 .extended_lut = "off";
defparam \ShiftLeft2~9 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~9 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~9 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[9]~q ),
	.datae(!\ShiftLeft2~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~9 .extended_lut = "off";
defparam \data_reg~9 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~9 .shared_arith = "off";

dffeas \data_reg[9] (
	.clk(clk_clk),
	.d(\data_reg~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[9]~q ),
	.prn(vcc));
defparam \data_reg[9] .is_wysiwyg = "true";
defparam \data_reg[9] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~10 (
	.dataa(!q_a_10),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_10_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~10 .extended_lut = "off";
defparam \ShiftLeft2~10 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~10 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~10 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[10]~q ),
	.datae(!\ShiftLeft2~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~10 .extended_lut = "off";
defparam \data_reg~10 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~10 .shared_arith = "off";

dffeas \data_reg[10] (
	.clk(clk_clk),
	.d(\data_reg~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[10]~q ),
	.prn(vcc));
defparam \data_reg[10] .is_wysiwyg = "true";
defparam \data_reg[10] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~11 (
	.dataa(!q_a_11),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_11_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~11 .extended_lut = "off";
defparam \ShiftLeft2~11 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~11 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~11 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[11]~q ),
	.datae(!\ShiftLeft2~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~11 .extended_lut = "off";
defparam \data_reg~11 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~11 .shared_arith = "off";

dffeas \data_reg[11] (
	.clk(clk_clk),
	.d(\data_reg~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[11]~q ),
	.prn(vcc));
defparam \data_reg[11] .is_wysiwyg = "true";
defparam \data_reg[11] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~12 (
	.dataa(!q_a_12),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_12_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~12 .extended_lut = "off";
defparam \ShiftLeft2~12 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~12 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~12 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[12]~q ),
	.datae(!\ShiftLeft2~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~12 .extended_lut = "off";
defparam \data_reg~12 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~12 .shared_arith = "off";

dffeas \data_reg[12] (
	.clk(clk_clk),
	.d(\data_reg~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[12]~q ),
	.prn(vcc));
defparam \data_reg[12] .is_wysiwyg = "true";
defparam \data_reg[12] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~13 (
	.dataa(!q_a_13),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_13_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~13 .extended_lut = "off";
defparam \ShiftLeft2~13 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~13 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~13 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[13]~q ),
	.datae(!\ShiftLeft2~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~13 .extended_lut = "off";
defparam \data_reg~13 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~13 .shared_arith = "off";

dffeas \data_reg[13] (
	.clk(clk_clk),
	.d(\data_reg~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[13]~q ),
	.prn(vcc));
defparam \data_reg[13] .is_wysiwyg = "true";
defparam \data_reg[13] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~14 (
	.dataa(!q_a_14),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_14_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~14 .extended_lut = "off";
defparam \ShiftLeft2~14 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~14 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~14 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[14]~q ),
	.datae(!\ShiftLeft2~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~14 .extended_lut = "off";
defparam \data_reg~14 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~14 .shared_arith = "off";

dffeas \data_reg[14] (
	.clk(clk_clk),
	.d(\data_reg~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[14]~q ),
	.prn(vcc));
defparam \data_reg[14] .is_wysiwyg = "true";
defparam \data_reg[14] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft2~15 (
	.dataa(!q_a_15),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!mem_15_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft2~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft2~15 .extended_lut = "off";
defparam \ShiftLeft2~15 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \ShiftLeft2~15 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~15 (
	.dataa(!source_addr_1),
	.datab(!source_addr_11),
	.datac(!mem_19_0),
	.datad(!\data_reg[15]~q ),
	.datae(!\ShiftLeft2~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~15 .extended_lut = "off";
defparam \data_reg~15 .lut_mask = 64'h00FFB8FF00FFB8FF;
defparam \data_reg~15 .shared_arith = "off";

dffeas \data_reg[15] (
	.clk(clk_clk),
	.d(\data_reg~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\always10~0_combout ),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(\data_reg[15]~q ),
	.prn(vcc));
defparam \data_reg[15] .is_wysiwyg = "true";
defparam \data_reg[15] .power_up = "low";

endmodule

module system_system_mm_interconnect_0_cmd_mux (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	Add4,
	Add5,
	Add41,
	Add51,
	Add42,
	Add52,
	Add43,
	Add53,
	Add44,
	Add54,
	src_data_66,
	saved_grant_1,
	saved_grant_0,
	src_data_78,
	src_data_79,
	src_data_77,
	in_ready,
	nxt_out_eop,
	nxt_out_eop1,
	nxt_in_ready,
	nxt_in_ready1,
	sink1_ready1,
	nxt_in_ready2,
	src_valid,
	write_addr_data_both_valid,
	r_sync_rst,
	WideOr11,
	src_payload,
	Add1,
	src_payload1,
	Add3,
	src_data_70,
	sop_enable,
	write_cp_data_69,
	src_payload2,
	src_data_69,
	burst_bytecount_5,
	Add6,
	Add2,
	src_data_68,
	burst_bytecount_4,
	Add61,
	Add21,
	src_data_67,
	burst_bytecount_3,
	Add22,
	burst_bytecount_2,
	src_data_65,
	src_payload3,
	src_payload4,
	src_payload5,
	Add11,
	src_payload6,
	Add31,
	src_data_71,
	src_payload7,
	LessThan12,
	src_payload8,
	src_data_72,
	address_burst_2,
	src_data_38,
	src_payload9,
	src_data_73,
	address_burst_3,
	src_data_39,
	src_payload10,
	src_payload11,
	src_data_74,
	src_payload12,
	src_payload_0,
	src_data_701,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_711,
	src_data_721,
	src_data_731,
	src_payload13,
	src_data_741,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	Add4;
input 	Add5;
input 	Add41;
input 	Add51;
input 	Add42;
input 	Add52;
input 	Add43;
input 	Add53;
input 	Add44;
input 	Add54;
output 	src_data_66;
output 	saved_grant_1;
output 	saved_grant_0;
output 	src_data_78;
output 	src_data_79;
output 	src_data_77;
input 	in_ready;
input 	nxt_out_eop;
input 	nxt_out_eop1;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	sink1_ready1;
input 	nxt_in_ready2;
output 	src_valid;
input 	write_addr_data_both_valid;
input 	r_sync_rst;
output 	WideOr11;
output 	src_payload;
input 	Add1;
output 	src_payload1;
input 	Add3;
output 	src_data_70;
input 	sop_enable;
input 	write_cp_data_69;
output 	src_payload2;
output 	src_data_69;
input 	burst_bytecount_5;
input 	Add6;
input 	Add2;
output 	src_data_68;
input 	burst_bytecount_4;
input 	Add61;
input 	Add21;
output 	src_data_67;
input 	burst_bytecount_3;
input 	Add22;
input 	burst_bytecount_2;
output 	src_data_65;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
input 	Add11;
output 	src_payload6;
input 	Add31;
output 	src_data_71;
output 	src_payload7;
input 	LessThan12;
output 	src_payload8;
output 	src_data_72;
input 	address_burst_2;
output 	src_data_38;
output 	src_payload9;
output 	src_data_73;
input 	address_burst_3;
output 	src_data_39;
output 	src_payload10;
output 	src_payload11;
output 	src_data_74;
output 	src_payload12;
output 	src_payload_0;
output 	src_data_701;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_711;
output 	src_data_721;
output 	src_data_731;
output 	src_payload13;
output 	src_data_741;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \always6~0_combout ;
wire \last_cycle~0_combout ;
wire \update_grant~0_combout ;
wire \src_payload~2_combout ;
wire \src_payload~1_combout ;
wire \src_payload~4_combout ;
wire \src_data[74]~0_combout ;
wire \src_data[70]~1_combout ;
wire \src_data[70]~2_combout ;
wire \src_data[71]~4_combout ;
wire \src_data[72]~6_combout ;
wire \src_data[72]~7_combout ;
wire \src_data[73]~9_combout ;
wire \src_data[73]~10_combout ;
wire \src_data[74]~12_combout ;
wire \src_payload~16_combout ;
wire \src_data[70]~14_combout ;
wire \src_data[71]~16_combout ;
wire \src_data[72]~18_combout ;
wire \src_data[73]~20_combout ;
wire \src_data[74]~22_combout ;


system_altera_merlin_arbitrator arb(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.in_ready(in_ready),
	.nxt_in_ready(nxt_in_ready1),
	.nxt_in_ready1(nxt_in_ready2),
	.write_addr_data_both_valid(write_addr_data_both_valid),
	.grant_1(\arb|grant[1]~0_combout ),
	.reset(r_sync_rst),
	.always6(\always6~0_combout ),
	.last_cycle(\last_cycle~0_combout ),
	.grant_0(\arb|grant[0]~1_combout ),
	.clk(clk_clk));

cyclonev_lcell_comb \src_data[66]~24 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!Add22),
	.datac(!burst_bytecount_3),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!saved_grant_1),
	.datag(!h2f_lw_AWLEN_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[66]~24 .extended_lut = "on";
defparam \src_data[66]~24 .lut_mask = 64'h005A000F337B333F;
defparam \src_data[66]~24 .shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb sink1_ready(
	.dataa(!saved_grant_1),
	.datab(!in_ready),
	.datac(!nxt_out_eop),
	.datad(!nxt_out_eop1),
	.datae(!nxt_in_ready),
	.dataf(!nxt_in_ready1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink1_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam sink1_ready.extended_lut = "off";
defparam sink1_ready.lut_mask = 64'h4444444400000444;
defparam sink1_ready.shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!saved_grant_1),
	.datae(!saved_grant_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h0055035700550357;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h0202020202020202;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!\src_payload~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h0080008000800080;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~3 (
	.dataa(!Add5),
	.datab(!\src_payload~1_combout ),
	.datac(!src_payload1),
	.datad(!\src_payload~4_combout ),
	.datae(!\src_data[70]~1_combout ),
	.dataf(!\src_data[70]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~3 .extended_lut = "off";
defparam \src_data[70]~3 .lut_mask = 64'hEE0E000000000000;
defparam \src_data[70]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h0000000100000001;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[69] (
	.dataa(!saved_grant_0),
	.datab(!write_cp_data_69),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[69] .extended_lut = "off";
defparam \src_data[69] .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \src_data[69] .shared_arith = "off";

cyclonev_lcell_comb \src_data[68] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!sop_enable),
	.datad(!burst_bytecount_5),
	.datae(!Add6),
	.dataf(!Add2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[68] .extended_lut = "off";
defparam \src_data[68] .lut_mask = 64'h0003303355577577;
defparam \src_data[68] .shared_arith = "off";

cyclonev_lcell_comb \src_data[67] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!sop_enable),
	.datad(!burst_bytecount_4),
	.datae(!Add61),
	.dataf(!Add21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[67] .extended_lut = "off";
defparam \src_data[67] .lut_mask = 64'h0003303355577577;
defparam \src_data[67] .shared_arith = "off";

cyclonev_lcell_comb \src_data[65] (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_AWLEN_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!burst_bytecount_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_65),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[65] .extended_lut = "off";
defparam \src_data[65] .lut_mask = 64'h0ACE0A0A0ACE0AFF;
defparam \src_data[65] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h0606060606060606;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h000001FE000001FE;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add41),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h0202020202020202;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!Add11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h8000800080008000;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~5 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~4_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add51),
	.datae(!src_payload6),
	.dataf(!\src_data[71]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~5 .extended_lut = "off";
defparam \src_data[71]~5 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[71]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add42),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h0202020202020202;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!LessThan12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h8000800080008000;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~8 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~4_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add52),
	.datae(!src_payload8),
	.dataf(!\src_data[72]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~8 .extended_lut = "off";
defparam \src_data[72]~8 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[72]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!h2f_lw_AWADDR_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!address_burst_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h05370505053705FF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add43),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h0202020202020202;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~11 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_data[70]~2_combout ),
	.datac(!Add53),
	.datad(!\src_data[73]~9_combout ),
	.datae(!\src_data[73]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~11 .extended_lut = "off";
defparam \src_data[73]~11 .lut_mask = 64'hC8000000C8000000;
defparam \src_data[73]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!h2f_lw_AWADDR_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!address_burst_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h05370505053705FF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add44),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h0202020202020202;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!\src_payload~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h80E880E880E880E8;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~13 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~4_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add54),
	.datae(!src_payload11),
	.dataf(!\src_data[74]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~13 .extended_lut = "off";
defparam \src_data[74]~13 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[74]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_ARADDR_4),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~15 (
	.dataa(!Add5),
	.datab(!\src_payload~1_combout ),
	.datac(!Add4),
	.datad(!\src_payload~16_combout ),
	.datae(!\src_data[70]~1_combout ),
	.dataf(!\src_data[70]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_701),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~15 .extended_lut = "off";
defparam \src_data[70]~15 .lut_mask = 64'hFFFFFFFF111FFFFF;
defparam \src_data[70]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0537053705370537;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0537053705370537;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0537053705370537;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~17 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~16_combout ),
	.datac(!Add51),
	.datad(!Add41),
	.datae(!\src_data[71]~4_combout ),
	.dataf(!\src_data[71]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_711),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~17 .extended_lut = "off";
defparam \src_data[71]~17 .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[71]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~19 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~16_combout ),
	.datac(!Add52),
	.datad(!Add42),
	.datae(!\src_data[72]~7_combout ),
	.dataf(!\src_data[72]~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_721),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~19 .extended_lut = "off";
defparam \src_data[72]~19 .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[72]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~21 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~16_combout ),
	.datac(!Add53),
	.datad(!Add43),
	.datae(!\src_data[73]~10_combout ),
	.dataf(!\src_data[73]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_731),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~21 .extended_lut = "off";
defparam \src_data[73]~21 .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[73]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h8080808080808080;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~23 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~16_combout ),
	.datac(!Add54),
	.datad(!Add44),
	.datae(!\src_data[74]~12_combout ),
	.dataf(!\src_data[74]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_741),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~23 .extended_lut = "off";
defparam \src_data[74]~23 .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[74]~23 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \always6~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!saved_grant_1),
	.datae(!saved_grant_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hFFAAFCA800000000;
defparam \always6~0 .shared_arith = "off";

cyclonev_lcell_comb \last_cycle~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WLAST_0),
	.datad(!h2f_lw_WVALID_0),
	.datae(!saved_grant_1),
	.dataf(!saved_grant_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_cycle~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~0 .extended_lut = "off";
defparam \last_cycle~0 .lut_mask = 64'h0000555500035577;
defparam \last_cycle~0 .shared_arith = "off";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready2),
	.datac(!nxt_in_ready1),
	.datad(!\always6~0_combout ),
	.datae(!\last_cycle~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'h00FFA2FF00FFA2FF;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(!h2f_lw_AWSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h80FF0F0030004000;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h2222222222222222;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~0 .extended_lut = "off";
defparam \src_data[74]~0 .lut_mask = 64'h80FF0F0030004000;
defparam \src_data[74]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~1 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!h2f_lw_ARLEN_3),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!saved_grant_1),
	.datae(!Add3),
	.dataf(!\src_data[74]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~1 .extended_lut = "off";
defparam \src_data[70]~1 .lut_mask = 64'h0055005500150055;
defparam \src_data[70]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~2 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_AWBURST_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~2 .extended_lut = "off";
defparam \src_data[70]~2 .lut_mask = 64'h0537053705370537;
defparam \src_data[70]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~4 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!h2f_lw_ARLEN_3),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!saved_grant_1),
	.datae(!Add3),
	.dataf(!Add31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[71]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~4 .extended_lut = "off";
defparam \src_data[71]~4 .lut_mask = 64'h0015005500550055;
defparam \src_data[71]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~6 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~6 .extended_lut = "off";
defparam \src_data[72]~6 .lut_mask = 64'h0F003000400080FF;
defparam \src_data[72]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~7 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!h2f_lw_ARLEN_3),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!saved_grant_1),
	.datae(!Add3),
	.dataf(!\src_data[72]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~7 .extended_lut = "off";
defparam \src_data[72]~7 .lut_mask = 64'h0015005500550055;
defparam \src_data[72]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~9 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!h2f_lw_ARLEN_3),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!saved_grant_1),
	.datae(!Add3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~9 .extended_lut = "off";
defparam \src_data[73]~9 .lut_mask = 64'h0015005500150055;
defparam \src_data[73]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~10 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!h2f_lw_AWLEN_3),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!saved_grant_0),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~10 .extended_lut = "off";
defparam \src_data[73]~10 .lut_mask = 64'h0015005500150055;
defparam \src_data[73]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~12 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!h2f_lw_ARLEN_3),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!saved_grant_1),
	.datae(!Add3),
	.dataf(!\src_data[74]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~12 .extended_lut = "off";
defparam \src_data[74]~12 .lut_mask = 64'h0015005500010015;
defparam \src_data[74]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h2222222222222222;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~14 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!\src_payload~2_combout ),
	.datae(!\src_payload~4_combout ),
	.dataf(!\src_data[70]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~14 .extended_lut = "off";
defparam \src_data[70]~14 .lut_mask = 64'hFFFF008000000000;
defparam \src_data[70]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~16 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!Add11),
	.datae(!\src_payload~4_combout ),
	.dataf(!\src_data[70]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[71]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~16 .extended_lut = "off";
defparam \src_data[71]~16 .lut_mask = 64'hFFFF800000000000;
defparam \src_data[71]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~18 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!\src_payload~4_combout ),
	.datae(!\src_data[70]~2_combout ),
	.dataf(!LessThan12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~18 .extended_lut = "off";
defparam \src_data[72]~18 .lut_mask = 64'hFF800000FF000000;
defparam \src_data[72]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~20 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!h2f_lw_ARLEN_3),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!saved_grant_1),
	.datae(!Add3),
	.dataf(!\src_data[70]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~20 .extended_lut = "off";
defparam \src_data[73]~20 .lut_mask = 64'hFFEAFFAA00000000;
defparam \src_data[73]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~22 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!Add1),
	.datad(!\src_payload~2_combout ),
	.datae(!\src_payload~4_combout ),
	.dataf(!\src_data[70]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~22 .extended_lut = "off";
defparam \src_data[74]~22 .lut_mask = 64'hFFFF80E800000000;
defparam \src_data[74]~22 .shared_arith = "off";

endmodule

module system_altera_merlin_arbitrator (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	in_ready,
	nxt_in_ready,
	nxt_in_ready1,
	write_addr_data_both_valid,
	grant_1,
	reset,
	always6,
	last_cycle,
	grant_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
input 	in_ready;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	write_addr_data_both_valid;
output 	grant_1;
input 	reset;
input 	always6;
input 	last_cycle;
output 	grant_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!write_addr_data_both_valid),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h4505450545054505;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!write_addr_data_both_valid),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h3302330233023302;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hA8A8A8A8A8A8A8A8;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!always6),
	.datae(!last_cycle),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h00FFA2FF00000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module system_system_mm_interconnect_0_rsp_demux (
	always10,
	out_valid,
	mem_95_0,
	mem_39_0,
	last_packet_beat,
	mem_41_0,
	src0_valid,
	src0_valid1,
	src1_valid)/* synthesis synthesis_greybox=0 */;
input 	always10;
input 	out_valid;
input 	mem_95_0;
input 	mem_39_0;
input 	last_packet_beat;
input 	mem_41_0;
output 	src0_valid;
output 	src0_valid1;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!mem_39_0),
	.datab(!mem_41_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h2222222222222222;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~1 (
	.dataa(!out_valid),
	.datab(!mem_95_0),
	.datac(!last_packet_beat),
	.datad(!always10),
	.datae(!src0_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~1 .extended_lut = "off";
defparam \src0_valid~1 .lut_mask = 64'h000020AA000020AA;
defparam \src0_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!out_valid),
	.datab(!mem_95_0),
	.datac(!last_packet_beat),
	.datad(!always10),
	.datae(!src0_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h20AA000020AA0000;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module system_system_pll_0 (
	outclk_wire_1,
	outclk_wire_0,
	merged_reset,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_1;
output 	outclk_wire_0;
input 	merged_reset;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altera_pll_1 altera_pll_i(
	.outclk({outclk_wire_1,outclk_wire_0}),
	.rst(merged_reset),
	.refclk(clk_clk));

endmodule

module system_altera_pll_1 (
	outclk,
	rst,
	refclk)/* synthesis synthesis_greybox=0 */;
output 	[1:0] outclk;
input 	rst;
input 	refclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fboutclk_wire[0] ;


generic_pll \general[1].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[1]),
	.fboutclk(),
	.locked(),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[1].gpll .clock_name_global = "false";
defparam \general[1].gpll .duty_cycle = 50;
defparam \general[1].gpll .fractional_vco_multiplier = "false";
defparam \general[1].gpll .output_clock_frequency = "108.0 mhz";
defparam \general[1].gpll .phase_shift = "8796 ps";
defparam \general[1].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[1].gpll .simulation_type = "timing";

generic_pll \general[0].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[0]),
	.fboutclk(\fboutclk_wire[0] ),
	.locked(),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[0].gpll .clock_name_global = "false";
defparam \general[0].gpll .duty_cycle = 50;
defparam \general[0].gpll .fractional_vco_multiplier = "false";
defparam \general[0].gpll .output_clock_frequency = "108.0 mhz";
defparam \general[0].gpll .phase_shift = "0 ps";
defparam \general[0].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[0].gpll .simulation_type = "timing";

endmodule

module system_system_ram (
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	q_a_8,
	q_b_8,
	q_a_9,
	q_b_9,
	q_a_10,
	q_b_10,
	q_a_11,
	q_b_11,
	q_a_12,
	q_b_12,
	q_a_13,
	q_b_13,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	in_data_reg_0,
	int_nxt_addr_reg_dly_1,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	m0_write,
	r_early_rst,
	source0_data_16,
	source0_data_17,
	clk_clk,
	ram_conduit_chipselect,
	ram_conduit_write,
	ram_conduit_clken,
	ram_conduit_writedata_0,
	ram_conduit_address_0,
	ram_conduit_address_1,
	ram_conduit_address_2,
	ram_conduit_address_3,
	ram_conduit_byteenable_0,
	ram_conduit_writedata_1,
	ram_conduit_writedata_2,
	ram_conduit_writedata_3,
	ram_conduit_writedata_4,
	ram_conduit_writedata_5,
	ram_conduit_writedata_6,
	ram_conduit_writedata_7,
	ram_conduit_writedata_8,
	ram_conduit_byteenable_1,
	ram_conduit_writedata_9,
	ram_conduit_writedata_10,
	ram_conduit_writedata_11,
	ram_conduit_writedata_12,
	ram_conduit_writedata_13,
	ram_conduit_writedata_14,
	ram_conduit_writedata_15)/* synthesis synthesis_greybox=0 */;
output 	q_a_0;
output 	q_b_0;
output 	q_a_1;
output 	q_b_1;
output 	q_a_2;
output 	q_b_2;
output 	q_a_3;
output 	q_b_3;
output 	q_a_4;
output 	q_b_4;
output 	q_a_5;
output 	q_b_5;
output 	q_a_6;
output 	q_b_6;
output 	q_a_7;
output 	q_b_7;
output 	q_a_8;
output 	q_b_8;
output 	q_a_9;
output 	q_b_9;
output 	q_a_10;
output 	q_b_10;
output 	q_a_11;
output 	q_b_11;
output 	q_a_12;
output 	q_b_12;
output 	q_a_13;
output 	q_b_13;
output 	q_a_14;
output 	q_b_14;
output 	q_a_15;
output 	q_b_15;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_1;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_4;
input 	in_data_reg_1;
input 	in_data_reg_2;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	m0_write;
input 	r_early_rst;
input 	source0_data_16;
input 	source0_data_17;
input 	clk_clk;
input 	ram_conduit_chipselect;
input 	ram_conduit_write;
input 	ram_conduit_clken;
input 	ram_conduit_writedata_0;
input 	ram_conduit_address_0;
input 	ram_conduit_address_1;
input 	ram_conduit_address_2;
input 	ram_conduit_address_3;
input 	ram_conduit_byteenable_0;
input 	ram_conduit_writedata_1;
input 	ram_conduit_writedata_2;
input 	ram_conduit_writedata_3;
input 	ram_conduit_writedata_4;
input 	ram_conduit_writedata_5;
input 	ram_conduit_writedata_6;
input 	ram_conduit_writedata_7;
input 	ram_conduit_writedata_8;
input 	ram_conduit_byteenable_1;
input 	ram_conduit_writedata_9;
input 	ram_conduit_writedata_10;
input 	ram_conduit_writedata_11;
input 	ram_conduit_writedata_12;
input 	ram_conduit_writedata_13;
input 	ram_conduit_writedata_14;
input 	ram_conduit_writedata_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren2~combout ;
wire \clocken1~combout ;


system_altsyncram_1 the_altsyncram(
	.q_a({q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({in_data_reg_15,in_data_reg_14,in_data_reg_13,in_data_reg_12,in_data_reg_11,in_data_reg_10,in_data_reg_9,in_data_reg_8,in_data_reg_7,in_data_reg_6,in_data_reg_5,in_data_reg_4,in_data_reg_3,in_data_reg_2,in_data_reg_1,in_data_reg_0}),
	.address_a({int_nxt_addr_reg_dly_4,int_nxt_addr_reg_dly_3,int_nxt_addr_reg_dly_2,int_nxt_addr_reg_dly_1}),
	.wren_a(m0_write),
	.wren_b(\wren2~combout ),
	.clocken0(r_early_rst),
	.clocken1(\clocken1~combout ),
	.byteena_a({source0_data_17,source0_data_16}),
	.clock0(clk_clk),
	.data_b({ram_conduit_writedata_15,ram_conduit_writedata_14,ram_conduit_writedata_13,ram_conduit_writedata_12,ram_conduit_writedata_11,ram_conduit_writedata_10,ram_conduit_writedata_9,ram_conduit_writedata_8,ram_conduit_writedata_7,ram_conduit_writedata_6,
ram_conduit_writedata_5,ram_conduit_writedata_4,ram_conduit_writedata_3,ram_conduit_writedata_2,ram_conduit_writedata_1,ram_conduit_writedata_0}),
	.address_b({ram_conduit_address_3,ram_conduit_address_2,ram_conduit_address_1,ram_conduit_address_0}),
	.byteena_b({ram_conduit_byteenable_1,ram_conduit_byteenable_0}));

cyclonev_lcell_comb wren2(
	.dataa(!ram_conduit_chipselect),
	.datab(!ram_conduit_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren2~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wren2.extended_lut = "off";
defparam wren2.lut_mask = 64'h1111111111111111;
defparam wren2.shared_arith = "off";

cyclonev_lcell_comb clocken1(
	.dataa(!r_early_rst),
	.datab(!ram_conduit_clken),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clocken1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam clocken1.extended_lut = "off";
defparam clocken1.lut_mask = 64'h2222222222222222;
defparam clocken1.shared_arith = "off";

endmodule

module system_altsyncram_1 (
	q_a,
	q_b,
	data_a,
	address_a,
	wren_a,
	wren_b,
	clocken0,
	clocken1,
	byteena_a,
	clock0,
	data_b,
	address_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
output 	[15:0] q_a;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	wren_b;
input 	clocken0;
input 	clocken1;
input 	[1:0] byteena_a;
input 	clock0;
input 	[15:0] data_b;
input 	[3:0] address_b;
input 	[1:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



system_altsyncram_2v72 auto_generated(
	.q_a({q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.wren_b(wren_b),
	.clocken0(clocken0),
	.clocken1(clocken1),
	.byteena_a({byteena_a[1],byteena_a[0]}),
	.clock0(clock0),
	.clock1(clock0),
	.data_b({data_b[15],data_b[14],data_b[13],data_b[12],data_b[11],data_b[10],data_b[9],data_b[8],data_b[7],data_b[6],data_b[5],data_b[4],data_b[3],data_b[2],data_b[1],data_b[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.byteena_b({byteena_b[1],byteena_b[0]}));

endmodule

module system_altsyncram_2v72 (
	q_a,
	q_b,
	data_a,
	address_a,
	wren_a,
	wren_b,
	clocken0,
	clocken1,
	byteena_a,
	clock0,
	clock1,
	data_b,
	address_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
output 	[15:0] q_a;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	wren_b;
input 	clocken0;
input 	clocken1;
input 	[1:0] byteena_a;
input 	clock0;
input 	clock1;
input 	[15:0] data_b;
input 	[3:0] address_b;
input 	[1:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "system_ram.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_byte_enable_clock = "clock1";
defparam ram_block1a0.port_b_byte_enable_mask_width = 1;
defparam ram_block1a0.port_b_byte_size = 1;
defparam ram_block1a0.port_b_data_in_clock = "clock1";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.port_b_write_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "0000";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "system_ram.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_byte_enable_clock = "clock1";
defparam ram_block1a1.port_b_byte_enable_mask_width = 1;
defparam ram_block1a1.port_b_byte_size = 1;
defparam ram_block1a1.port_b_data_in_clock = "clock1";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.port_b_write_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "0000";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "system_ram.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_byte_enable_clock = "clock1";
defparam ram_block1a2.port_b_byte_enable_mask_width = 1;
defparam ram_block1a2.port_b_byte_size = 1;
defparam ram_block1a2.port_b_data_in_clock = "clock1";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.port_b_write_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "0000";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "system_ram.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_byte_enable_clock = "clock1";
defparam ram_block1a3.port_b_byte_enable_mask_width = 1;
defparam ram_block1a3.port_b_byte_size = 1;
defparam ram_block1a3.port_b_data_in_clock = "clock1";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.port_b_write_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "0000";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "system_ram.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_byte_enable_clock = "clock1";
defparam ram_block1a4.port_b_byte_enable_mask_width = 1;
defparam ram_block1a4.port_b_byte_size = 1;
defparam ram_block1a4.port_b_data_in_clock = "clock1";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.port_b_write_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "0000";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "system_ram.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_byte_enable_clock = "clock1";
defparam ram_block1a5.port_b_byte_enable_mask_width = 1;
defparam ram_block1a5.port_b_byte_size = 1;
defparam ram_block1a5.port_b_data_in_clock = "clock1";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.port_b_write_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "0000";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "system_ram.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_byte_enable_clock = "clock1";
defparam ram_block1a6.port_b_byte_enable_mask_width = 1;
defparam ram_block1a6.port_b_byte_size = 1;
defparam ram_block1a6.port_b_data_in_clock = "clock1";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.port_b_write_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "0000";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "system_ram.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_byte_enable_clock = "clock1";
defparam ram_block1a7.port_b_byte_enable_mask_width = 1;
defparam ram_block1a7.port_b_byte_size = 1;
defparam ram_block1a7.port_b_data_in_clock = "clock1";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.port_b_write_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "0000";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "system_ram.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_byte_enable_clock = "clock1";
defparam ram_block1a8.port_b_byte_enable_mask_width = 1;
defparam ram_block1a8.port_b_byte_size = 1;
defparam ram_block1a8.port_b_data_in_clock = "clock1";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.port_b_write_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "0000";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "system_ram.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_byte_enable_clock = "clock1";
defparam ram_block1a9.port_b_byte_enable_mask_width = 1;
defparam ram_block1a9.port_b_byte_size = 1;
defparam ram_block1a9.port_b_data_in_clock = "clock1";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.port_b_write_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "0000";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "system_ram.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_byte_enable_clock = "clock1";
defparam ram_block1a10.port_b_byte_enable_mask_width = 1;
defparam ram_block1a10.port_b_byte_size = 1;
defparam ram_block1a10.port_b_data_in_clock = "clock1";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.port_b_write_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "0000";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "system_ram.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_byte_enable_clock = "clock1";
defparam ram_block1a11.port_b_byte_enable_mask_width = 1;
defparam ram_block1a11.port_b_byte_size = 1;
defparam ram_block1a11.port_b_data_in_clock = "clock1";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.port_b_write_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "0000";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "system_ram.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_byte_enable_clock = "clock1";
defparam ram_block1a12.port_b_byte_enable_mask_width = 1;
defparam ram_block1a12.port_b_byte_size = 1;
defparam ram_block1a12.port_b_data_in_clock = "clock1";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.port_b_write_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "0000";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "system_ram.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_byte_enable_clock = "clock1";
defparam ram_block1a13.port_b_byte_enable_mask_width = 1;
defparam ram_block1a13.port_b_byte_size = 1;
defparam ram_block1a13.port_b_data_in_clock = "clock1";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.port_b_write_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "0000";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "system_ram.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_byte_enable_clock = "clock1";
defparam ram_block1a14.port_b_byte_enable_mask_width = 1;
defparam ram_block1a14.port_b_byte_size = 1;
defparam ram_block1a14.port_b_data_in_clock = "clock1";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.port_b_write_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "0000";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "system_ram.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "system_ram:ram|altsyncram:the_altsyncram|altsyncram_2v72:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_byte_enable_clock = "clock1";
defparam ram_block1a15.port_b_byte_enable_mask_width = 1;
defparam ram_block1a15.port_b_byte_size = 1;
defparam ram_block1a15.port_b_data_in_clock = "clock1";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.port_b_write_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "0000";

endmodule
