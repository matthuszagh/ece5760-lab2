/* top.v
 *
 * A top level module to instantiate the other submodules and control their operation.
 */

module top (
            // Clocks
            input CLOCK_50,

            )
