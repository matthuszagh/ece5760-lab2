
module system (
	clk_clk,
	reset_reset_n,
	vga_clk_ext_clk,
	vga_clk_int_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		vga_clk_ext_clk;
	output		vga_clk_int_clk;
endmodule
